
`include "sample_manager.sv"
`include "csv_file_dump.sv"
`include "df_fifo_monitor.sv"
`include "df_process_monitor.sv"
`include "nodf_module_monitor.sv"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_MPSQ.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_MPSQ.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_MPSQ.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_makeSuperPoint_alignedToLine_2_fu_23088.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_makeSuperPoint_alignedToLine_2_fu_23088.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_makeSuperPoint_alignedToLine_2_fu_23088.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_makeSuperPoint_alignedToLine_2_fu_23088.grp_mSP_findBounds_fu_21923.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_makeSuperPoint_alignedToLine_2_fu_23088.grp_mSP_findBounds_fu_21923.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_makeSuperPoint_alignedToLine_2_fu_23088.grp_mSP_findBounds_fu_21923.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = 1'b0;
    assign module_intf_9.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_add_patch_patches_parameters_fu_8850.ap_ready;
    assign module_intf_9.ap_done = 1'b0;
    assign module_intf_9.ap_continue = 1'b0;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = 1'b0;
    assign module_intf_10.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8914.ap_ready;
    assign module_intf_10.ap_done = 1'b0;
    assign module_intf_10.ap_continue = 1'b0;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = 1'b0;
    assign module_intf_11.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8921.ap_ready;
    assign module_intf_11.ap_done = 1'b0;
    assign module_intf_11.ap_continue = 1'b0;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = 1'b0;
    assign module_intf_12.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8928.ap_ready;
    assign module_intf_12.ap_done = 1'b0;
    assign module_intf_12.ap_continue = 1'b0;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = 1'b0;
    assign module_intf_13.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8935.ap_ready;
    assign module_intf_13.ap_done = 1'b0;
    assign module_intf_13.ap_continue = 1'b0;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = 1'b0;
    assign module_intf_14.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8942.ap_ready;
    assign module_intf_14.ap_done = 1'b0;
    assign module_intf_14.ap_continue = 1'b0;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = 1'b0;
    assign module_intf_15.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8949.ap_ready;
    assign module_intf_15.ap_done = 1'b0;
    assign module_intf_15.ap_continue = 1'b0;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = 1'b0;
    assign module_intf_16.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8956.ap_ready;
    assign module_intf_16.ap_done = 1'b0;
    assign module_intf_16.ap_continue = 1'b0;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = 1'b0;
    assign module_intf_17.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8963.ap_ready;
    assign module_intf_17.ap_done = 1'b0;
    assign module_intf_17.ap_continue = 1'b0;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = 1'b0;
    assign module_intf_18.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8970.ap_ready;
    assign module_intf_18.ap_done = 1'b0;
    assign module_intf_18.ap_continue = 1'b0;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = 1'b0;
    assign module_intf_19.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8977.ap_ready;
    assign module_intf_19.ap_done = 1'b0;
    assign module_intf_19.ap_continue = 1'b0;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = 1'b0;
    assign module_intf_20.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8984.ap_ready;
    assign module_intf_20.ap_done = 1'b0;
    assign module_intf_20.ap_continue = 1'b0;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = 1'b0;
    assign module_intf_21.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8991.ap_ready;
    assign module_intf_21.ap_done = 1'b0;
    assign module_intf_21.ap_continue = 1'b0;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = 1'b0;
    assign module_intf_22.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8998.ap_ready;
    assign module_intf_22.ap_done = 1'b0;
    assign module_intf_22.ap_continue = 1'b0;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = 1'b0;
    assign module_intf_23.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9005.ap_ready;
    assign module_intf_23.ap_done = 1'b0;
    assign module_intf_23.ap_continue = 1'b0;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = 1'b0;
    assign module_intf_24.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9012.ap_ready;
    assign module_intf_24.ap_done = 1'b0;
    assign module_intf_24.ap_continue = 1'b0;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = 1'b0;
    assign module_intf_25.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9019.ap_ready;
    assign module_intf_25.ap_done = 1'b0;
    assign module_intf_25.ap_continue = 1'b0;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = 1'b0;
    assign module_intf_26.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9026.ap_ready;
    assign module_intf_26.ap_done = 1'b0;
    assign module_intf_26.ap_continue = 1'b0;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = 1'b0;
    assign module_intf_27.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9033.ap_ready;
    assign module_intf_27.ap_done = 1'b0;
    assign module_intf_27.ap_continue = 1'b0;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = 1'b0;
    assign module_intf_28.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9040.ap_ready;
    assign module_intf_28.ap_done = 1'b0;
    assign module_intf_28.ap_continue = 1'b0;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = 1'b0;
    assign module_intf_29.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9047.ap_ready;
    assign module_intf_29.ap_done = 1'b0;
    assign module_intf_29.ap_continue = 1'b0;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = 1'b0;
    assign module_intf_30.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9054.ap_ready;
    assign module_intf_30.ap_done = 1'b0;
    assign module_intf_30.ap_continue = 1'b0;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = 1'b0;
    assign module_intf_31.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9061.ap_ready;
    assign module_intf_31.ap_done = 1'b0;
    assign module_intf_31.ap_continue = 1'b0;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = 1'b0;
    assign module_intf_32.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9068.ap_ready;
    assign module_intf_32.ap_done = 1'b0;
    assign module_intf_32.ap_continue = 1'b0;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = 1'b0;
    assign module_intf_33.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9075.ap_ready;
    assign module_intf_33.ap_done = 1'b0;
    assign module_intf_33.ap_continue = 1'b0;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = 1'b0;
    assign module_intf_34.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9082.ap_ready;
    assign module_intf_34.ap_done = 1'b0;
    assign module_intf_34.ap_continue = 1'b0;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = 1'b0;
    assign module_intf_35.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9089.ap_ready;
    assign module_intf_35.ap_done = 1'b0;
    assign module_intf_35.ap_continue = 1'b0;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = 1'b0;
    assign module_intf_36.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9096.ap_ready;
    assign module_intf_36.ap_done = 1'b0;
    assign module_intf_36.ap_continue = 1'b0;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = 1'b0;
    assign module_intf_37.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9103.ap_ready;
    assign module_intf_37.ap_done = 1'b0;
    assign module_intf_37.ap_continue = 1'b0;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = 1'b0;
    assign module_intf_38.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9110.ap_ready;
    assign module_intf_38.ap_done = 1'b0;
    assign module_intf_38.ap_continue = 1'b0;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = 1'b0;
    assign module_intf_39.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9117.ap_ready;
    assign module_intf_39.ap_done = 1'b0;
    assign module_intf_39.ap_continue = 1'b0;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = 1'b0;
    assign module_intf_40.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9124.ap_ready;
    assign module_intf_40.ap_done = 1'b0;
    assign module_intf_40.ap_continue = 1'b0;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = 1'b0;
    assign module_intf_41.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9131.ap_ready;
    assign module_intf_41.ap_done = 1'b0;
    assign module_intf_41.ap_continue = 1'b0;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = 1'b0;
    assign module_intf_42.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9138.ap_ready;
    assign module_intf_42.ap_done = 1'b0;
    assign module_intf_42.ap_continue = 1'b0;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = 1'b0;
    assign module_intf_43.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9145.ap_ready;
    assign module_intf_43.ap_done = 1'b0;
    assign module_intf_43.ap_continue = 1'b0;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = 1'b0;
    assign module_intf_44.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9152.ap_ready;
    assign module_intf_44.ap_done = 1'b0;
    assign module_intf_44.ap_continue = 1'b0;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = 1'b0;
    assign module_intf_45.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9159.ap_ready;
    assign module_intf_45.ap_done = 1'b0;
    assign module_intf_45.ap_continue = 1'b0;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = 1'b0;
    assign module_intf_46.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9166.ap_ready;
    assign module_intf_46.ap_done = 1'b0;
    assign module_intf_46.ap_continue = 1'b0;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = 1'b0;
    assign module_intf_47.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9173.ap_ready;
    assign module_intf_47.ap_done = 1'b0;
    assign module_intf_47.ap_continue = 1'b0;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = 1'b0;
    assign module_intf_48.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9180.ap_ready;
    assign module_intf_48.ap_done = 1'b0;
    assign module_intf_48.ap_continue = 1'b0;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = 1'b0;
    assign module_intf_49.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9187.ap_ready;
    assign module_intf_49.ap_done = 1'b0;
    assign module_intf_49.ap_continue = 1'b0;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = 1'b0;
    assign module_intf_50.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9194.ap_ready;
    assign module_intf_50.ap_done = 1'b0;
    assign module_intf_50.ap_continue = 1'b0;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = 1'b0;
    assign module_intf_51.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9201.ap_ready;
    assign module_intf_51.ap_done = 1'b0;
    assign module_intf_51.ap_continue = 1'b0;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = 1'b0;
    assign module_intf_52.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9208.ap_ready;
    assign module_intf_52.ap_done = 1'b0;
    assign module_intf_52.ap_continue = 1'b0;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = 1'b0;
    assign module_intf_53.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9215.ap_ready;
    assign module_intf_53.ap_done = 1'b0;
    assign module_intf_53.ap_continue = 1'b0;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = 1'b0;
    assign module_intf_54.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9222.ap_ready;
    assign module_intf_54.ap_done = 1'b0;
    assign module_intf_54.ap_continue = 1'b0;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = 1'b0;
    assign module_intf_55.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9229.ap_ready;
    assign module_intf_55.ap_done = 1'b0;
    assign module_intf_55.ap_continue = 1'b0;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = 1'b0;
    assign module_intf_56.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9236.ap_ready;
    assign module_intf_56.ap_done = 1'b0;
    assign module_intf_56.ap_continue = 1'b0;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = 1'b0;
    assign module_intf_57.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9243.ap_ready;
    assign module_intf_57.ap_done = 1'b0;
    assign module_intf_57.ap_continue = 1'b0;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;
    nodf_module_intf module_intf_58(clock,reset);
    assign module_intf_58.ap_start = 1'b0;
    assign module_intf_58.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9250.ap_ready;
    assign module_intf_58.ap_done = 1'b0;
    assign module_intf_58.ap_continue = 1'b0;
    assign module_intf_58.finish = finish;
    csv_file_dump mstatus_csv_dumper_58;
    nodf_module_monitor module_monitor_58;
    nodf_module_intf module_intf_59(clock,reset);
    assign module_intf_59.ap_start = 1'b0;
    assign module_intf_59.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9257.ap_ready;
    assign module_intf_59.ap_done = 1'b0;
    assign module_intf_59.ap_continue = 1'b0;
    assign module_intf_59.finish = finish;
    csv_file_dump mstatus_csv_dumper_59;
    nodf_module_monitor module_monitor_59;
    nodf_module_intf module_intf_60(clock,reset);
    assign module_intf_60.ap_start = 1'b0;
    assign module_intf_60.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9264.ap_ready;
    assign module_intf_60.ap_done = 1'b0;
    assign module_intf_60.ap_continue = 1'b0;
    assign module_intf_60.finish = finish;
    csv_file_dump mstatus_csv_dumper_60;
    nodf_module_monitor module_monitor_60;
    nodf_module_intf module_intf_61(clock,reset);
    assign module_intf_61.ap_start = 1'b0;
    assign module_intf_61.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9271.ap_ready;
    assign module_intf_61.ap_done = 1'b0;
    assign module_intf_61.ap_continue = 1'b0;
    assign module_intf_61.finish = finish;
    csv_file_dump mstatus_csv_dumper_61;
    nodf_module_monitor module_monitor_61;
    nodf_module_intf module_intf_62(clock,reset);
    assign module_intf_62.ap_start = 1'b0;
    assign module_intf_62.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9278.ap_ready;
    assign module_intf_62.ap_done = 1'b0;
    assign module_intf_62.ap_continue = 1'b0;
    assign module_intf_62.finish = finish;
    csv_file_dump mstatus_csv_dumper_62;
    nodf_module_monitor module_monitor_62;
    nodf_module_intf module_intf_63(clock,reset);
    assign module_intf_63.ap_start = 1'b0;
    assign module_intf_63.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9285.ap_ready;
    assign module_intf_63.ap_done = 1'b0;
    assign module_intf_63.ap_continue = 1'b0;
    assign module_intf_63.finish = finish;
    csv_file_dump mstatus_csv_dumper_63;
    nodf_module_monitor module_monitor_63;
    nodf_module_intf module_intf_64(clock,reset);
    assign module_intf_64.ap_start = 1'b0;
    assign module_intf_64.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9292.ap_ready;
    assign module_intf_64.ap_done = 1'b0;
    assign module_intf_64.ap_continue = 1'b0;
    assign module_intf_64.finish = finish;
    csv_file_dump mstatus_csv_dumper_64;
    nodf_module_monitor module_monitor_64;
    nodf_module_intf module_intf_65(clock,reset);
    assign module_intf_65.ap_start = 1'b0;
    assign module_intf_65.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9299.ap_ready;
    assign module_intf_65.ap_done = 1'b0;
    assign module_intf_65.ap_continue = 1'b0;
    assign module_intf_65.finish = finish;
    csv_file_dump mstatus_csv_dumper_65;
    nodf_module_monitor module_monitor_65;
    nodf_module_intf module_intf_66(clock,reset);
    assign module_intf_66.ap_start = 1'b0;
    assign module_intf_66.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9306.ap_ready;
    assign module_intf_66.ap_done = 1'b0;
    assign module_intf_66.ap_continue = 1'b0;
    assign module_intf_66.finish = finish;
    csv_file_dump mstatus_csv_dumper_66;
    nodf_module_monitor module_monitor_66;
    nodf_module_intf module_intf_67(clock,reset);
    assign module_intf_67.ap_start = 1'b0;
    assign module_intf_67.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9313.ap_ready;
    assign module_intf_67.ap_done = 1'b0;
    assign module_intf_67.ap_continue = 1'b0;
    assign module_intf_67.finish = finish;
    csv_file_dump mstatus_csv_dumper_67;
    nodf_module_monitor module_monitor_67;
    nodf_module_intf module_intf_68(clock,reset);
    assign module_intf_68.ap_start = 1'b0;
    assign module_intf_68.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9320.ap_ready;
    assign module_intf_68.ap_done = 1'b0;
    assign module_intf_68.ap_continue = 1'b0;
    assign module_intf_68.finish = finish;
    csv_file_dump mstatus_csv_dumper_68;
    nodf_module_monitor module_monitor_68;
    nodf_module_intf module_intf_69(clock,reset);
    assign module_intf_69.ap_start = 1'b0;
    assign module_intf_69.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9327.ap_ready;
    assign module_intf_69.ap_done = 1'b0;
    assign module_intf_69.ap_continue = 1'b0;
    assign module_intf_69.finish = finish;
    csv_file_dump mstatus_csv_dumper_69;
    nodf_module_monitor module_monitor_69;
    nodf_module_intf module_intf_70(clock,reset);
    assign module_intf_70.ap_start = 1'b0;
    assign module_intf_70.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9334.ap_ready;
    assign module_intf_70.ap_done = 1'b0;
    assign module_intf_70.ap_continue = 1'b0;
    assign module_intf_70.finish = finish;
    csv_file_dump mstatus_csv_dumper_70;
    nodf_module_monitor module_monitor_70;
    nodf_module_intf module_intf_71(clock,reset);
    assign module_intf_71.ap_start = 1'b0;
    assign module_intf_71.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9341.ap_ready;
    assign module_intf_71.ap_done = 1'b0;
    assign module_intf_71.ap_continue = 1'b0;
    assign module_intf_71.finish = finish;
    csv_file_dump mstatus_csv_dumper_71;
    nodf_module_monitor module_monitor_71;
    nodf_module_intf module_intf_72(clock,reset);
    assign module_intf_72.ap_start = 1'b0;
    assign module_intf_72.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9348.ap_ready;
    assign module_intf_72.ap_done = 1'b0;
    assign module_intf_72.ap_continue = 1'b0;
    assign module_intf_72.finish = finish;
    csv_file_dump mstatus_csv_dumper_72;
    nodf_module_monitor module_monitor_72;
    nodf_module_intf module_intf_73(clock,reset);
    assign module_intf_73.ap_start = 1'b0;
    assign module_intf_73.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9355.ap_ready;
    assign module_intf_73.ap_done = 1'b0;
    assign module_intf_73.ap_continue = 1'b0;
    assign module_intf_73.finish = finish;
    csv_file_dump mstatus_csv_dumper_73;
    nodf_module_monitor module_monitor_73;
    nodf_module_intf module_intf_74(clock,reset);
    assign module_intf_74.ap_start = 1'b0;
    assign module_intf_74.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9362.ap_ready;
    assign module_intf_74.ap_done = 1'b0;
    assign module_intf_74.ap_continue = 1'b0;
    assign module_intf_74.finish = finish;
    csv_file_dump mstatus_csv_dumper_74;
    nodf_module_monitor module_monitor_74;
    nodf_module_intf module_intf_75(clock,reset);
    assign module_intf_75.ap_start = 1'b0;
    assign module_intf_75.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9369.ap_ready;
    assign module_intf_75.ap_done = 1'b0;
    assign module_intf_75.ap_continue = 1'b0;
    assign module_intf_75.finish = finish;
    csv_file_dump mstatus_csv_dumper_75;
    nodf_module_monitor module_monitor_75;
    nodf_module_intf module_intf_76(clock,reset);
    assign module_intf_76.ap_start = 1'b0;
    assign module_intf_76.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9376.ap_ready;
    assign module_intf_76.ap_done = 1'b0;
    assign module_intf_76.ap_continue = 1'b0;
    assign module_intf_76.finish = finish;
    csv_file_dump mstatus_csv_dumper_76;
    nodf_module_monitor module_monitor_76;
    nodf_module_intf module_intf_77(clock,reset);
    assign module_intf_77.ap_start = 1'b0;
    assign module_intf_77.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9383.ap_ready;
    assign module_intf_77.ap_done = 1'b0;
    assign module_intf_77.ap_continue = 1'b0;
    assign module_intf_77.finish = finish;
    csv_file_dump mstatus_csv_dumper_77;
    nodf_module_monitor module_monitor_77;
    nodf_module_intf module_intf_78(clock,reset);
    assign module_intf_78.ap_start = 1'b0;
    assign module_intf_78.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9390.ap_ready;
    assign module_intf_78.ap_done = 1'b0;
    assign module_intf_78.ap_continue = 1'b0;
    assign module_intf_78.finish = finish;
    csv_file_dump mstatus_csv_dumper_78;
    nodf_module_monitor module_monitor_78;
    nodf_module_intf module_intf_79(clock,reset);
    assign module_intf_79.ap_start = 1'b0;
    assign module_intf_79.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9397.ap_ready;
    assign module_intf_79.ap_done = 1'b0;
    assign module_intf_79.ap_continue = 1'b0;
    assign module_intf_79.finish = finish;
    csv_file_dump mstatus_csv_dumper_79;
    nodf_module_monitor module_monitor_79;
    nodf_module_intf module_intf_80(clock,reset);
    assign module_intf_80.ap_start = 1'b0;
    assign module_intf_80.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9404.ap_ready;
    assign module_intf_80.ap_done = 1'b0;
    assign module_intf_80.ap_continue = 1'b0;
    assign module_intf_80.finish = finish;
    csv_file_dump mstatus_csv_dumper_80;
    nodf_module_monitor module_monitor_80;
    nodf_module_intf module_intf_81(clock,reset);
    assign module_intf_81.ap_start = 1'b0;
    assign module_intf_81.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9411.ap_ready;
    assign module_intf_81.ap_done = 1'b0;
    assign module_intf_81.ap_continue = 1'b0;
    assign module_intf_81.finish = finish;
    csv_file_dump mstatus_csv_dumper_81;
    nodf_module_monitor module_monitor_81;
    nodf_module_intf module_intf_82(clock,reset);
    assign module_intf_82.ap_start = 1'b0;
    assign module_intf_82.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9418.ap_ready;
    assign module_intf_82.ap_done = 1'b0;
    assign module_intf_82.ap_continue = 1'b0;
    assign module_intf_82.finish = finish;
    csv_file_dump mstatus_csv_dumper_82;
    nodf_module_monitor module_monitor_82;
    nodf_module_intf module_intf_83(clock,reset);
    assign module_intf_83.ap_start = 1'b0;
    assign module_intf_83.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9425.ap_ready;
    assign module_intf_83.ap_done = 1'b0;
    assign module_intf_83.ap_continue = 1'b0;
    assign module_intf_83.finish = finish;
    csv_file_dump mstatus_csv_dumper_83;
    nodf_module_monitor module_monitor_83;
    nodf_module_intf module_intf_84(clock,reset);
    assign module_intf_84.ap_start = 1'b0;
    assign module_intf_84.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9432.ap_ready;
    assign module_intf_84.ap_done = 1'b0;
    assign module_intf_84.ap_continue = 1'b0;
    assign module_intf_84.finish = finish;
    csv_file_dump mstatus_csv_dumper_84;
    nodf_module_monitor module_monitor_84;
    nodf_module_intf module_intf_85(clock,reset);
    assign module_intf_85.ap_start = 1'b0;
    assign module_intf_85.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9439.ap_ready;
    assign module_intf_85.ap_done = 1'b0;
    assign module_intf_85.ap_continue = 1'b0;
    assign module_intf_85.finish = finish;
    csv_file_dump mstatus_csv_dumper_85;
    nodf_module_monitor module_monitor_85;
    nodf_module_intf module_intf_86(clock,reset);
    assign module_intf_86.ap_start = 1'b0;
    assign module_intf_86.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9446.ap_ready;
    assign module_intf_86.ap_done = 1'b0;
    assign module_intf_86.ap_continue = 1'b0;
    assign module_intf_86.finish = finish;
    csv_file_dump mstatus_csv_dumper_86;
    nodf_module_monitor module_monitor_86;
    nodf_module_intf module_intf_87(clock,reset);
    assign module_intf_87.ap_start = 1'b0;
    assign module_intf_87.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9453.ap_ready;
    assign module_intf_87.ap_done = 1'b0;
    assign module_intf_87.ap_continue = 1'b0;
    assign module_intf_87.finish = finish;
    csv_file_dump mstatus_csv_dumper_87;
    nodf_module_monitor module_monitor_87;
    nodf_module_intf module_intf_88(clock,reset);
    assign module_intf_88.ap_start = 1'b0;
    assign module_intf_88.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9460.ap_ready;
    assign module_intf_88.ap_done = 1'b0;
    assign module_intf_88.ap_continue = 1'b0;
    assign module_intf_88.finish = finish;
    csv_file_dump mstatus_csv_dumper_88;
    nodf_module_monitor module_monitor_88;
    nodf_module_intf module_intf_89(clock,reset);
    assign module_intf_89.ap_start = 1'b0;
    assign module_intf_89.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9467.ap_ready;
    assign module_intf_89.ap_done = 1'b0;
    assign module_intf_89.ap_continue = 1'b0;
    assign module_intf_89.finish = finish;
    csv_file_dump mstatus_csv_dumper_89;
    nodf_module_monitor module_monitor_89;
    nodf_module_intf module_intf_90(clock,reset);
    assign module_intf_90.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.ap_start;
    assign module_intf_90.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.ap_ready;
    assign module_intf_90.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.ap_done;
    assign module_intf_90.ap_continue = 1'b1;
    assign module_intf_90.finish = finish;
    csv_file_dump mstatus_csv_dumper_90;
    nodf_module_monitor module_monitor_90;
    nodf_module_intf module_intf_91(clock,reset);
    assign module_intf_91.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_start;
    assign module_intf_91.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_ready;
    assign module_intf_91.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_done;
    assign module_intf_91.ap_continue = 1'b1;
    assign module_intf_91.finish = finish;
    csv_file_dump mstatus_csv_dumper_91;
    nodf_module_monitor module_monitor_91;
    nodf_module_intf module_intf_92(clock,reset);
    assign module_intf_92.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_start;
    assign module_intf_92.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_ready;
    assign module_intf_92.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_done;
    assign module_intf_92.ap_continue = 1'b1;
    assign module_intf_92.finish = finish;
    csv_file_dump mstatus_csv_dumper_92;
    nodf_module_monitor module_monitor_92;
    nodf_module_intf module_intf_93(clock,reset);
    assign module_intf_93.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_start;
    assign module_intf_93.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_ready;
    assign module_intf_93.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_done;
    assign module_intf_93.ap_continue = 1'b1;
    assign module_intf_93.finish = finish;
    csv_file_dump mstatus_csv_dumper_93;
    nodf_module_monitor module_monitor_93;
    nodf_module_intf module_intf_94(clock,reset);
    assign module_intf_94.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_start;
    assign module_intf_94.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_ready;
    assign module_intf_94.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_done;
    assign module_intf_94.ap_continue = 1'b1;
    assign module_intf_94.finish = finish;
    csv_file_dump mstatus_csv_dumper_94;
    nodf_module_monitor module_monitor_94;
    nodf_module_intf module_intf_95(clock,reset);
    assign module_intf_95.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_start;
    assign module_intf_95.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_ready;
    assign module_intf_95.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_makePatch_alignedToLine_2_fu_30135.grp_wedgePatch_init_fu_29542.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_done;
    assign module_intf_95.ap_continue = 1'b1;
    assign module_intf_95.finish = finish;
    csv_file_dump mstatus_csv_dumper_95;
    nodf_module_monitor module_monitor_95;
    nodf_module_intf module_intf_96(clock,reset);
    assign module_intf_96.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_delete_patch_fu_33340.ap_start;
    assign module_intf_96.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_delete_patch_fu_33340.ap_ready;
    assign module_intf_96.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_delete_patch_fu_33340.ap_done;
    assign module_intf_96.ap_continue = 1'b1;
    assign module_intf_96.finish = finish;
    csv_file_dump mstatus_csv_dumper_96;
    nodf_module_monitor module_monitor_96;
    nodf_module_intf module_intf_97(clock,reset);
    assign module_intf_97.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_delete_patch_fu_33340.grp_delete_patch_patches_parameters_fu_10118.ap_start;
    assign module_intf_97.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_delete_patch_fu_33340.grp_delete_patch_patches_parameters_fu_10118.ap_ready;
    assign module_intf_97.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_delete_patch_fu_33340.grp_delete_patch_patches_parameters_fu_10118.ap_done;
    assign module_intf_97.ap_continue = 1'b1;
    assign module_intf_97.finish = finish;
    csv_file_dump mstatus_csv_dumper_97;
    nodf_module_monitor module_monitor_97;
    nodf_module_intf module_intf_98(clock,reset);
    assign module_intf_98.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_get_index_from_z_fu_33740.ap_start;
    assign module_intf_98.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_get_index_from_z_fu_33740.ap_ready;
    assign module_intf_98.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_solveComplmentaryPatch_fu_36470.grp_get_index_from_z_fu_33740.ap_done;
    assign module_intf_98.ap_continue = 1'b1;
    assign module_intf_98.finish = finish;
    csv_file_dump mstatus_csv_dumper_98;
    nodf_module_monitor module_monitor_98;
    nodf_module_intf module_intf_99(clock,reset);
    assign module_intf_99.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.ap_start;
    assign module_intf_99.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.ap_ready;
    assign module_intf_99.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.ap_done;
    assign module_intf_99.ap_continue = 1'b1;
    assign module_intf_99.finish = finish;
    csv_file_dump mstatus_csv_dumper_99;
    nodf_module_monitor module_monitor_99;
    nodf_module_intf module_intf_100(clock,reset);
    assign module_intf_100.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.ap_start;
    assign module_intf_100.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.ap_ready;
    assign module_intf_100.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.ap_done;
    assign module_intf_100.ap_continue = 1'b1;
    assign module_intf_100.finish = finish;
    csv_file_dump mstatus_csv_dumper_100;
    nodf_module_monitor module_monitor_100;
    nodf_module_intf module_intf_101(clock,reset);
    assign module_intf_101.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_makeSuperPoint_alignedToLine_1_fu_23098.ap_start;
    assign module_intf_101.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_makeSuperPoint_alignedToLine_1_fu_23098.ap_ready;
    assign module_intf_101.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_makeSuperPoint_alignedToLine_1_fu_23098.ap_done;
    assign module_intf_101.ap_continue = 1'b1;
    assign module_intf_101.finish = finish;
    csv_file_dump mstatus_csv_dumper_101;
    nodf_module_monitor module_monitor_101;
    nodf_module_intf module_intf_102(clock,reset);
    assign module_intf_102.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_makeSuperPoint_alignedToLine_1_fu_23098.grp_mSP_findBounds_fu_21935.ap_start;
    assign module_intf_102.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_makeSuperPoint_alignedToLine_1_fu_23098.grp_mSP_findBounds_fu_21935.ap_ready;
    assign module_intf_102.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_makeSuperPoint_alignedToLine_1_fu_23098.grp_mSP_findBounds_fu_21935.ap_done;
    assign module_intf_102.ap_continue = 1'b1;
    assign module_intf_102.finish = finish;
    csv_file_dump mstatus_csv_dumper_102;
    nodf_module_monitor module_monitor_102;
    nodf_module_intf module_intf_103(clock,reset);
    assign module_intf_103.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.ap_start;
    assign module_intf_103.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.ap_ready;
    assign module_intf_103.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.ap_done;
    assign module_intf_103.ap_continue = 1'b1;
    assign module_intf_103.finish = finish;
    csv_file_dump mstatus_csv_dumper_103;
    nodf_module_monitor module_monitor_103;
    nodf_module_intf module_intf_104(clock,reset);
    assign module_intf_104.ap_start = 1'b0;
    assign module_intf_104.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_add_patch_patches_parameters_fu_8850.ap_ready;
    assign module_intf_104.ap_done = 1'b0;
    assign module_intf_104.ap_continue = 1'b0;
    assign module_intf_104.finish = finish;
    csv_file_dump mstatus_csv_dumper_104;
    nodf_module_monitor module_monitor_104;
    nodf_module_intf module_intf_105(clock,reset);
    assign module_intf_105.ap_start = 1'b0;
    assign module_intf_105.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8914.ap_ready;
    assign module_intf_105.ap_done = 1'b0;
    assign module_intf_105.ap_continue = 1'b0;
    assign module_intf_105.finish = finish;
    csv_file_dump mstatus_csv_dumper_105;
    nodf_module_monitor module_monitor_105;
    nodf_module_intf module_intf_106(clock,reset);
    assign module_intf_106.ap_start = 1'b0;
    assign module_intf_106.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8921.ap_ready;
    assign module_intf_106.ap_done = 1'b0;
    assign module_intf_106.ap_continue = 1'b0;
    assign module_intf_106.finish = finish;
    csv_file_dump mstatus_csv_dumper_106;
    nodf_module_monitor module_monitor_106;
    nodf_module_intf module_intf_107(clock,reset);
    assign module_intf_107.ap_start = 1'b0;
    assign module_intf_107.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8928.ap_ready;
    assign module_intf_107.ap_done = 1'b0;
    assign module_intf_107.ap_continue = 1'b0;
    assign module_intf_107.finish = finish;
    csv_file_dump mstatus_csv_dumper_107;
    nodf_module_monitor module_monitor_107;
    nodf_module_intf module_intf_108(clock,reset);
    assign module_intf_108.ap_start = 1'b0;
    assign module_intf_108.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8935.ap_ready;
    assign module_intf_108.ap_done = 1'b0;
    assign module_intf_108.ap_continue = 1'b0;
    assign module_intf_108.finish = finish;
    csv_file_dump mstatus_csv_dumper_108;
    nodf_module_monitor module_monitor_108;
    nodf_module_intf module_intf_109(clock,reset);
    assign module_intf_109.ap_start = 1'b0;
    assign module_intf_109.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8942.ap_ready;
    assign module_intf_109.ap_done = 1'b0;
    assign module_intf_109.ap_continue = 1'b0;
    assign module_intf_109.finish = finish;
    csv_file_dump mstatus_csv_dumper_109;
    nodf_module_monitor module_monitor_109;
    nodf_module_intf module_intf_110(clock,reset);
    assign module_intf_110.ap_start = 1'b0;
    assign module_intf_110.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8949.ap_ready;
    assign module_intf_110.ap_done = 1'b0;
    assign module_intf_110.ap_continue = 1'b0;
    assign module_intf_110.finish = finish;
    csv_file_dump mstatus_csv_dumper_110;
    nodf_module_monitor module_monitor_110;
    nodf_module_intf module_intf_111(clock,reset);
    assign module_intf_111.ap_start = 1'b0;
    assign module_intf_111.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8956.ap_ready;
    assign module_intf_111.ap_done = 1'b0;
    assign module_intf_111.ap_continue = 1'b0;
    assign module_intf_111.finish = finish;
    csv_file_dump mstatus_csv_dumper_111;
    nodf_module_monitor module_monitor_111;
    nodf_module_intf module_intf_112(clock,reset);
    assign module_intf_112.ap_start = 1'b0;
    assign module_intf_112.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8963.ap_ready;
    assign module_intf_112.ap_done = 1'b0;
    assign module_intf_112.ap_continue = 1'b0;
    assign module_intf_112.finish = finish;
    csv_file_dump mstatus_csv_dumper_112;
    nodf_module_monitor module_monitor_112;
    nodf_module_intf module_intf_113(clock,reset);
    assign module_intf_113.ap_start = 1'b0;
    assign module_intf_113.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8970.ap_ready;
    assign module_intf_113.ap_done = 1'b0;
    assign module_intf_113.ap_continue = 1'b0;
    assign module_intf_113.finish = finish;
    csv_file_dump mstatus_csv_dumper_113;
    nodf_module_monitor module_monitor_113;
    nodf_module_intf module_intf_114(clock,reset);
    assign module_intf_114.ap_start = 1'b0;
    assign module_intf_114.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8977.ap_ready;
    assign module_intf_114.ap_done = 1'b0;
    assign module_intf_114.ap_continue = 1'b0;
    assign module_intf_114.finish = finish;
    csv_file_dump mstatus_csv_dumper_114;
    nodf_module_monitor module_monitor_114;
    nodf_module_intf module_intf_115(clock,reset);
    assign module_intf_115.ap_start = 1'b0;
    assign module_intf_115.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8984.ap_ready;
    assign module_intf_115.ap_done = 1'b0;
    assign module_intf_115.ap_continue = 1'b0;
    assign module_intf_115.finish = finish;
    csv_file_dump mstatus_csv_dumper_115;
    nodf_module_monitor module_monitor_115;
    nodf_module_intf module_intf_116(clock,reset);
    assign module_intf_116.ap_start = 1'b0;
    assign module_intf_116.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8991.ap_ready;
    assign module_intf_116.ap_done = 1'b0;
    assign module_intf_116.ap_continue = 1'b0;
    assign module_intf_116.finish = finish;
    csv_file_dump mstatus_csv_dumper_116;
    nodf_module_monitor module_monitor_116;
    nodf_module_intf module_intf_117(clock,reset);
    assign module_intf_117.ap_start = 1'b0;
    assign module_intf_117.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8998.ap_ready;
    assign module_intf_117.ap_done = 1'b0;
    assign module_intf_117.ap_continue = 1'b0;
    assign module_intf_117.finish = finish;
    csv_file_dump mstatus_csv_dumper_117;
    nodf_module_monitor module_monitor_117;
    nodf_module_intf module_intf_118(clock,reset);
    assign module_intf_118.ap_start = 1'b0;
    assign module_intf_118.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9005.ap_ready;
    assign module_intf_118.ap_done = 1'b0;
    assign module_intf_118.ap_continue = 1'b0;
    assign module_intf_118.finish = finish;
    csv_file_dump mstatus_csv_dumper_118;
    nodf_module_monitor module_monitor_118;
    nodf_module_intf module_intf_119(clock,reset);
    assign module_intf_119.ap_start = 1'b0;
    assign module_intf_119.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9012.ap_ready;
    assign module_intf_119.ap_done = 1'b0;
    assign module_intf_119.ap_continue = 1'b0;
    assign module_intf_119.finish = finish;
    csv_file_dump mstatus_csv_dumper_119;
    nodf_module_monitor module_monitor_119;
    nodf_module_intf module_intf_120(clock,reset);
    assign module_intf_120.ap_start = 1'b0;
    assign module_intf_120.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9019.ap_ready;
    assign module_intf_120.ap_done = 1'b0;
    assign module_intf_120.ap_continue = 1'b0;
    assign module_intf_120.finish = finish;
    csv_file_dump mstatus_csv_dumper_120;
    nodf_module_monitor module_monitor_120;
    nodf_module_intf module_intf_121(clock,reset);
    assign module_intf_121.ap_start = 1'b0;
    assign module_intf_121.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9026.ap_ready;
    assign module_intf_121.ap_done = 1'b0;
    assign module_intf_121.ap_continue = 1'b0;
    assign module_intf_121.finish = finish;
    csv_file_dump mstatus_csv_dumper_121;
    nodf_module_monitor module_monitor_121;
    nodf_module_intf module_intf_122(clock,reset);
    assign module_intf_122.ap_start = 1'b0;
    assign module_intf_122.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9033.ap_ready;
    assign module_intf_122.ap_done = 1'b0;
    assign module_intf_122.ap_continue = 1'b0;
    assign module_intf_122.finish = finish;
    csv_file_dump mstatus_csv_dumper_122;
    nodf_module_monitor module_monitor_122;
    nodf_module_intf module_intf_123(clock,reset);
    assign module_intf_123.ap_start = 1'b0;
    assign module_intf_123.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9040.ap_ready;
    assign module_intf_123.ap_done = 1'b0;
    assign module_intf_123.ap_continue = 1'b0;
    assign module_intf_123.finish = finish;
    csv_file_dump mstatus_csv_dumper_123;
    nodf_module_monitor module_monitor_123;
    nodf_module_intf module_intf_124(clock,reset);
    assign module_intf_124.ap_start = 1'b0;
    assign module_intf_124.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9047.ap_ready;
    assign module_intf_124.ap_done = 1'b0;
    assign module_intf_124.ap_continue = 1'b0;
    assign module_intf_124.finish = finish;
    csv_file_dump mstatus_csv_dumper_124;
    nodf_module_monitor module_monitor_124;
    nodf_module_intf module_intf_125(clock,reset);
    assign module_intf_125.ap_start = 1'b0;
    assign module_intf_125.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9054.ap_ready;
    assign module_intf_125.ap_done = 1'b0;
    assign module_intf_125.ap_continue = 1'b0;
    assign module_intf_125.finish = finish;
    csv_file_dump mstatus_csv_dumper_125;
    nodf_module_monitor module_monitor_125;
    nodf_module_intf module_intf_126(clock,reset);
    assign module_intf_126.ap_start = 1'b0;
    assign module_intf_126.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9061.ap_ready;
    assign module_intf_126.ap_done = 1'b0;
    assign module_intf_126.ap_continue = 1'b0;
    assign module_intf_126.finish = finish;
    csv_file_dump mstatus_csv_dumper_126;
    nodf_module_monitor module_monitor_126;
    nodf_module_intf module_intf_127(clock,reset);
    assign module_intf_127.ap_start = 1'b0;
    assign module_intf_127.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9068.ap_ready;
    assign module_intf_127.ap_done = 1'b0;
    assign module_intf_127.ap_continue = 1'b0;
    assign module_intf_127.finish = finish;
    csv_file_dump mstatus_csv_dumper_127;
    nodf_module_monitor module_monitor_127;
    nodf_module_intf module_intf_128(clock,reset);
    assign module_intf_128.ap_start = 1'b0;
    assign module_intf_128.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9075.ap_ready;
    assign module_intf_128.ap_done = 1'b0;
    assign module_intf_128.ap_continue = 1'b0;
    assign module_intf_128.finish = finish;
    csv_file_dump mstatus_csv_dumper_128;
    nodf_module_monitor module_monitor_128;
    nodf_module_intf module_intf_129(clock,reset);
    assign module_intf_129.ap_start = 1'b0;
    assign module_intf_129.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9082.ap_ready;
    assign module_intf_129.ap_done = 1'b0;
    assign module_intf_129.ap_continue = 1'b0;
    assign module_intf_129.finish = finish;
    csv_file_dump mstatus_csv_dumper_129;
    nodf_module_monitor module_monitor_129;
    nodf_module_intf module_intf_130(clock,reset);
    assign module_intf_130.ap_start = 1'b0;
    assign module_intf_130.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9089.ap_ready;
    assign module_intf_130.ap_done = 1'b0;
    assign module_intf_130.ap_continue = 1'b0;
    assign module_intf_130.finish = finish;
    csv_file_dump mstatus_csv_dumper_130;
    nodf_module_monitor module_monitor_130;
    nodf_module_intf module_intf_131(clock,reset);
    assign module_intf_131.ap_start = 1'b0;
    assign module_intf_131.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9096.ap_ready;
    assign module_intf_131.ap_done = 1'b0;
    assign module_intf_131.ap_continue = 1'b0;
    assign module_intf_131.finish = finish;
    csv_file_dump mstatus_csv_dumper_131;
    nodf_module_monitor module_monitor_131;
    nodf_module_intf module_intf_132(clock,reset);
    assign module_intf_132.ap_start = 1'b0;
    assign module_intf_132.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9103.ap_ready;
    assign module_intf_132.ap_done = 1'b0;
    assign module_intf_132.ap_continue = 1'b0;
    assign module_intf_132.finish = finish;
    csv_file_dump mstatus_csv_dumper_132;
    nodf_module_monitor module_monitor_132;
    nodf_module_intf module_intf_133(clock,reset);
    assign module_intf_133.ap_start = 1'b0;
    assign module_intf_133.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9110.ap_ready;
    assign module_intf_133.ap_done = 1'b0;
    assign module_intf_133.ap_continue = 1'b0;
    assign module_intf_133.finish = finish;
    csv_file_dump mstatus_csv_dumper_133;
    nodf_module_monitor module_monitor_133;
    nodf_module_intf module_intf_134(clock,reset);
    assign module_intf_134.ap_start = 1'b0;
    assign module_intf_134.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9117.ap_ready;
    assign module_intf_134.ap_done = 1'b0;
    assign module_intf_134.ap_continue = 1'b0;
    assign module_intf_134.finish = finish;
    csv_file_dump mstatus_csv_dumper_134;
    nodf_module_monitor module_monitor_134;
    nodf_module_intf module_intf_135(clock,reset);
    assign module_intf_135.ap_start = 1'b0;
    assign module_intf_135.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9124.ap_ready;
    assign module_intf_135.ap_done = 1'b0;
    assign module_intf_135.ap_continue = 1'b0;
    assign module_intf_135.finish = finish;
    csv_file_dump mstatus_csv_dumper_135;
    nodf_module_monitor module_monitor_135;
    nodf_module_intf module_intf_136(clock,reset);
    assign module_intf_136.ap_start = 1'b0;
    assign module_intf_136.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9131.ap_ready;
    assign module_intf_136.ap_done = 1'b0;
    assign module_intf_136.ap_continue = 1'b0;
    assign module_intf_136.finish = finish;
    csv_file_dump mstatus_csv_dumper_136;
    nodf_module_monitor module_monitor_136;
    nodf_module_intf module_intf_137(clock,reset);
    assign module_intf_137.ap_start = 1'b0;
    assign module_intf_137.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9138.ap_ready;
    assign module_intf_137.ap_done = 1'b0;
    assign module_intf_137.ap_continue = 1'b0;
    assign module_intf_137.finish = finish;
    csv_file_dump mstatus_csv_dumper_137;
    nodf_module_monitor module_monitor_137;
    nodf_module_intf module_intf_138(clock,reset);
    assign module_intf_138.ap_start = 1'b0;
    assign module_intf_138.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9145.ap_ready;
    assign module_intf_138.ap_done = 1'b0;
    assign module_intf_138.ap_continue = 1'b0;
    assign module_intf_138.finish = finish;
    csv_file_dump mstatus_csv_dumper_138;
    nodf_module_monitor module_monitor_138;
    nodf_module_intf module_intf_139(clock,reset);
    assign module_intf_139.ap_start = 1'b0;
    assign module_intf_139.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9152.ap_ready;
    assign module_intf_139.ap_done = 1'b0;
    assign module_intf_139.ap_continue = 1'b0;
    assign module_intf_139.finish = finish;
    csv_file_dump mstatus_csv_dumper_139;
    nodf_module_monitor module_monitor_139;
    nodf_module_intf module_intf_140(clock,reset);
    assign module_intf_140.ap_start = 1'b0;
    assign module_intf_140.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9159.ap_ready;
    assign module_intf_140.ap_done = 1'b0;
    assign module_intf_140.ap_continue = 1'b0;
    assign module_intf_140.finish = finish;
    csv_file_dump mstatus_csv_dumper_140;
    nodf_module_monitor module_monitor_140;
    nodf_module_intf module_intf_141(clock,reset);
    assign module_intf_141.ap_start = 1'b0;
    assign module_intf_141.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9166.ap_ready;
    assign module_intf_141.ap_done = 1'b0;
    assign module_intf_141.ap_continue = 1'b0;
    assign module_intf_141.finish = finish;
    csv_file_dump mstatus_csv_dumper_141;
    nodf_module_monitor module_monitor_141;
    nodf_module_intf module_intf_142(clock,reset);
    assign module_intf_142.ap_start = 1'b0;
    assign module_intf_142.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9173.ap_ready;
    assign module_intf_142.ap_done = 1'b0;
    assign module_intf_142.ap_continue = 1'b0;
    assign module_intf_142.finish = finish;
    csv_file_dump mstatus_csv_dumper_142;
    nodf_module_monitor module_monitor_142;
    nodf_module_intf module_intf_143(clock,reset);
    assign module_intf_143.ap_start = 1'b0;
    assign module_intf_143.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9180.ap_ready;
    assign module_intf_143.ap_done = 1'b0;
    assign module_intf_143.ap_continue = 1'b0;
    assign module_intf_143.finish = finish;
    csv_file_dump mstatus_csv_dumper_143;
    nodf_module_monitor module_monitor_143;
    nodf_module_intf module_intf_144(clock,reset);
    assign module_intf_144.ap_start = 1'b0;
    assign module_intf_144.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9187.ap_ready;
    assign module_intf_144.ap_done = 1'b0;
    assign module_intf_144.ap_continue = 1'b0;
    assign module_intf_144.finish = finish;
    csv_file_dump mstatus_csv_dumper_144;
    nodf_module_monitor module_monitor_144;
    nodf_module_intf module_intf_145(clock,reset);
    assign module_intf_145.ap_start = 1'b0;
    assign module_intf_145.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9194.ap_ready;
    assign module_intf_145.ap_done = 1'b0;
    assign module_intf_145.ap_continue = 1'b0;
    assign module_intf_145.finish = finish;
    csv_file_dump mstatus_csv_dumper_145;
    nodf_module_monitor module_monitor_145;
    nodf_module_intf module_intf_146(clock,reset);
    assign module_intf_146.ap_start = 1'b0;
    assign module_intf_146.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9201.ap_ready;
    assign module_intf_146.ap_done = 1'b0;
    assign module_intf_146.ap_continue = 1'b0;
    assign module_intf_146.finish = finish;
    csv_file_dump mstatus_csv_dumper_146;
    nodf_module_monitor module_monitor_146;
    nodf_module_intf module_intf_147(clock,reset);
    assign module_intf_147.ap_start = 1'b0;
    assign module_intf_147.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9208.ap_ready;
    assign module_intf_147.ap_done = 1'b0;
    assign module_intf_147.ap_continue = 1'b0;
    assign module_intf_147.finish = finish;
    csv_file_dump mstatus_csv_dumper_147;
    nodf_module_monitor module_monitor_147;
    nodf_module_intf module_intf_148(clock,reset);
    assign module_intf_148.ap_start = 1'b0;
    assign module_intf_148.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9215.ap_ready;
    assign module_intf_148.ap_done = 1'b0;
    assign module_intf_148.ap_continue = 1'b0;
    assign module_intf_148.finish = finish;
    csv_file_dump mstatus_csv_dumper_148;
    nodf_module_monitor module_monitor_148;
    nodf_module_intf module_intf_149(clock,reset);
    assign module_intf_149.ap_start = 1'b0;
    assign module_intf_149.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9222.ap_ready;
    assign module_intf_149.ap_done = 1'b0;
    assign module_intf_149.ap_continue = 1'b0;
    assign module_intf_149.finish = finish;
    csv_file_dump mstatus_csv_dumper_149;
    nodf_module_monitor module_monitor_149;
    nodf_module_intf module_intf_150(clock,reset);
    assign module_intf_150.ap_start = 1'b0;
    assign module_intf_150.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9229.ap_ready;
    assign module_intf_150.ap_done = 1'b0;
    assign module_intf_150.ap_continue = 1'b0;
    assign module_intf_150.finish = finish;
    csv_file_dump mstatus_csv_dumper_150;
    nodf_module_monitor module_monitor_150;
    nodf_module_intf module_intf_151(clock,reset);
    assign module_intf_151.ap_start = 1'b0;
    assign module_intf_151.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9236.ap_ready;
    assign module_intf_151.ap_done = 1'b0;
    assign module_intf_151.ap_continue = 1'b0;
    assign module_intf_151.finish = finish;
    csv_file_dump mstatus_csv_dumper_151;
    nodf_module_monitor module_monitor_151;
    nodf_module_intf module_intf_152(clock,reset);
    assign module_intf_152.ap_start = 1'b0;
    assign module_intf_152.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9243.ap_ready;
    assign module_intf_152.ap_done = 1'b0;
    assign module_intf_152.ap_continue = 1'b0;
    assign module_intf_152.finish = finish;
    csv_file_dump mstatus_csv_dumper_152;
    nodf_module_monitor module_monitor_152;
    nodf_module_intf module_intf_153(clock,reset);
    assign module_intf_153.ap_start = 1'b0;
    assign module_intf_153.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9250.ap_ready;
    assign module_intf_153.ap_done = 1'b0;
    assign module_intf_153.ap_continue = 1'b0;
    assign module_intf_153.finish = finish;
    csv_file_dump mstatus_csv_dumper_153;
    nodf_module_monitor module_monitor_153;
    nodf_module_intf module_intf_154(clock,reset);
    assign module_intf_154.ap_start = 1'b0;
    assign module_intf_154.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9257.ap_ready;
    assign module_intf_154.ap_done = 1'b0;
    assign module_intf_154.ap_continue = 1'b0;
    assign module_intf_154.finish = finish;
    csv_file_dump mstatus_csv_dumper_154;
    nodf_module_monitor module_monitor_154;
    nodf_module_intf module_intf_155(clock,reset);
    assign module_intf_155.ap_start = 1'b0;
    assign module_intf_155.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9264.ap_ready;
    assign module_intf_155.ap_done = 1'b0;
    assign module_intf_155.ap_continue = 1'b0;
    assign module_intf_155.finish = finish;
    csv_file_dump mstatus_csv_dumper_155;
    nodf_module_monitor module_monitor_155;
    nodf_module_intf module_intf_156(clock,reset);
    assign module_intf_156.ap_start = 1'b0;
    assign module_intf_156.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9271.ap_ready;
    assign module_intf_156.ap_done = 1'b0;
    assign module_intf_156.ap_continue = 1'b0;
    assign module_intf_156.finish = finish;
    csv_file_dump mstatus_csv_dumper_156;
    nodf_module_monitor module_monitor_156;
    nodf_module_intf module_intf_157(clock,reset);
    assign module_intf_157.ap_start = 1'b0;
    assign module_intf_157.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9278.ap_ready;
    assign module_intf_157.ap_done = 1'b0;
    assign module_intf_157.ap_continue = 1'b0;
    assign module_intf_157.finish = finish;
    csv_file_dump mstatus_csv_dumper_157;
    nodf_module_monitor module_monitor_157;
    nodf_module_intf module_intf_158(clock,reset);
    assign module_intf_158.ap_start = 1'b0;
    assign module_intf_158.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9285.ap_ready;
    assign module_intf_158.ap_done = 1'b0;
    assign module_intf_158.ap_continue = 1'b0;
    assign module_intf_158.finish = finish;
    csv_file_dump mstatus_csv_dumper_158;
    nodf_module_monitor module_monitor_158;
    nodf_module_intf module_intf_159(clock,reset);
    assign module_intf_159.ap_start = 1'b0;
    assign module_intf_159.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9292.ap_ready;
    assign module_intf_159.ap_done = 1'b0;
    assign module_intf_159.ap_continue = 1'b0;
    assign module_intf_159.finish = finish;
    csv_file_dump mstatus_csv_dumper_159;
    nodf_module_monitor module_monitor_159;
    nodf_module_intf module_intf_160(clock,reset);
    assign module_intf_160.ap_start = 1'b0;
    assign module_intf_160.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9299.ap_ready;
    assign module_intf_160.ap_done = 1'b0;
    assign module_intf_160.ap_continue = 1'b0;
    assign module_intf_160.finish = finish;
    csv_file_dump mstatus_csv_dumper_160;
    nodf_module_monitor module_monitor_160;
    nodf_module_intf module_intf_161(clock,reset);
    assign module_intf_161.ap_start = 1'b0;
    assign module_intf_161.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9306.ap_ready;
    assign module_intf_161.ap_done = 1'b0;
    assign module_intf_161.ap_continue = 1'b0;
    assign module_intf_161.finish = finish;
    csv_file_dump mstatus_csv_dumper_161;
    nodf_module_monitor module_monitor_161;
    nodf_module_intf module_intf_162(clock,reset);
    assign module_intf_162.ap_start = 1'b0;
    assign module_intf_162.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9313.ap_ready;
    assign module_intf_162.ap_done = 1'b0;
    assign module_intf_162.ap_continue = 1'b0;
    assign module_intf_162.finish = finish;
    csv_file_dump mstatus_csv_dumper_162;
    nodf_module_monitor module_monitor_162;
    nodf_module_intf module_intf_163(clock,reset);
    assign module_intf_163.ap_start = 1'b0;
    assign module_intf_163.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9320.ap_ready;
    assign module_intf_163.ap_done = 1'b0;
    assign module_intf_163.ap_continue = 1'b0;
    assign module_intf_163.finish = finish;
    csv_file_dump mstatus_csv_dumper_163;
    nodf_module_monitor module_monitor_163;
    nodf_module_intf module_intf_164(clock,reset);
    assign module_intf_164.ap_start = 1'b0;
    assign module_intf_164.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9327.ap_ready;
    assign module_intf_164.ap_done = 1'b0;
    assign module_intf_164.ap_continue = 1'b0;
    assign module_intf_164.finish = finish;
    csv_file_dump mstatus_csv_dumper_164;
    nodf_module_monitor module_monitor_164;
    nodf_module_intf module_intf_165(clock,reset);
    assign module_intf_165.ap_start = 1'b0;
    assign module_intf_165.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9334.ap_ready;
    assign module_intf_165.ap_done = 1'b0;
    assign module_intf_165.ap_continue = 1'b0;
    assign module_intf_165.finish = finish;
    csv_file_dump mstatus_csv_dumper_165;
    nodf_module_monitor module_monitor_165;
    nodf_module_intf module_intf_166(clock,reset);
    assign module_intf_166.ap_start = 1'b0;
    assign module_intf_166.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9341.ap_ready;
    assign module_intf_166.ap_done = 1'b0;
    assign module_intf_166.ap_continue = 1'b0;
    assign module_intf_166.finish = finish;
    csv_file_dump mstatus_csv_dumper_166;
    nodf_module_monitor module_monitor_166;
    nodf_module_intf module_intf_167(clock,reset);
    assign module_intf_167.ap_start = 1'b0;
    assign module_intf_167.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9348.ap_ready;
    assign module_intf_167.ap_done = 1'b0;
    assign module_intf_167.ap_continue = 1'b0;
    assign module_intf_167.finish = finish;
    csv_file_dump mstatus_csv_dumper_167;
    nodf_module_monitor module_monitor_167;
    nodf_module_intf module_intf_168(clock,reset);
    assign module_intf_168.ap_start = 1'b0;
    assign module_intf_168.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9355.ap_ready;
    assign module_intf_168.ap_done = 1'b0;
    assign module_intf_168.ap_continue = 1'b0;
    assign module_intf_168.finish = finish;
    csv_file_dump mstatus_csv_dumper_168;
    nodf_module_monitor module_monitor_168;
    nodf_module_intf module_intf_169(clock,reset);
    assign module_intf_169.ap_start = 1'b0;
    assign module_intf_169.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9362.ap_ready;
    assign module_intf_169.ap_done = 1'b0;
    assign module_intf_169.ap_continue = 1'b0;
    assign module_intf_169.finish = finish;
    csv_file_dump mstatus_csv_dumper_169;
    nodf_module_monitor module_monitor_169;
    nodf_module_intf module_intf_170(clock,reset);
    assign module_intf_170.ap_start = 1'b0;
    assign module_intf_170.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9369.ap_ready;
    assign module_intf_170.ap_done = 1'b0;
    assign module_intf_170.ap_continue = 1'b0;
    assign module_intf_170.finish = finish;
    csv_file_dump mstatus_csv_dumper_170;
    nodf_module_monitor module_monitor_170;
    nodf_module_intf module_intf_171(clock,reset);
    assign module_intf_171.ap_start = 1'b0;
    assign module_intf_171.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9376.ap_ready;
    assign module_intf_171.ap_done = 1'b0;
    assign module_intf_171.ap_continue = 1'b0;
    assign module_intf_171.finish = finish;
    csv_file_dump mstatus_csv_dumper_171;
    nodf_module_monitor module_monitor_171;
    nodf_module_intf module_intf_172(clock,reset);
    assign module_intf_172.ap_start = 1'b0;
    assign module_intf_172.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9383.ap_ready;
    assign module_intf_172.ap_done = 1'b0;
    assign module_intf_172.ap_continue = 1'b0;
    assign module_intf_172.finish = finish;
    csv_file_dump mstatus_csv_dumper_172;
    nodf_module_monitor module_monitor_172;
    nodf_module_intf module_intf_173(clock,reset);
    assign module_intf_173.ap_start = 1'b0;
    assign module_intf_173.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9390.ap_ready;
    assign module_intf_173.ap_done = 1'b0;
    assign module_intf_173.ap_continue = 1'b0;
    assign module_intf_173.finish = finish;
    csv_file_dump mstatus_csv_dumper_173;
    nodf_module_monitor module_monitor_173;
    nodf_module_intf module_intf_174(clock,reset);
    assign module_intf_174.ap_start = 1'b0;
    assign module_intf_174.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9397.ap_ready;
    assign module_intf_174.ap_done = 1'b0;
    assign module_intf_174.ap_continue = 1'b0;
    assign module_intf_174.finish = finish;
    csv_file_dump mstatus_csv_dumper_174;
    nodf_module_monitor module_monitor_174;
    nodf_module_intf module_intf_175(clock,reset);
    assign module_intf_175.ap_start = 1'b0;
    assign module_intf_175.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9404.ap_ready;
    assign module_intf_175.ap_done = 1'b0;
    assign module_intf_175.ap_continue = 1'b0;
    assign module_intf_175.finish = finish;
    csv_file_dump mstatus_csv_dumper_175;
    nodf_module_monitor module_monitor_175;
    nodf_module_intf module_intf_176(clock,reset);
    assign module_intf_176.ap_start = 1'b0;
    assign module_intf_176.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9411.ap_ready;
    assign module_intf_176.ap_done = 1'b0;
    assign module_intf_176.ap_continue = 1'b0;
    assign module_intf_176.finish = finish;
    csv_file_dump mstatus_csv_dumper_176;
    nodf_module_monitor module_monitor_176;
    nodf_module_intf module_intf_177(clock,reset);
    assign module_intf_177.ap_start = 1'b0;
    assign module_intf_177.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9418.ap_ready;
    assign module_intf_177.ap_done = 1'b0;
    assign module_intf_177.ap_continue = 1'b0;
    assign module_intf_177.finish = finish;
    csv_file_dump mstatus_csv_dumper_177;
    nodf_module_monitor module_monitor_177;
    nodf_module_intf module_intf_178(clock,reset);
    assign module_intf_178.ap_start = 1'b0;
    assign module_intf_178.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9425.ap_ready;
    assign module_intf_178.ap_done = 1'b0;
    assign module_intf_178.ap_continue = 1'b0;
    assign module_intf_178.finish = finish;
    csv_file_dump mstatus_csv_dumper_178;
    nodf_module_monitor module_monitor_178;
    nodf_module_intf module_intf_179(clock,reset);
    assign module_intf_179.ap_start = 1'b0;
    assign module_intf_179.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9432.ap_ready;
    assign module_intf_179.ap_done = 1'b0;
    assign module_intf_179.ap_continue = 1'b0;
    assign module_intf_179.finish = finish;
    csv_file_dump mstatus_csv_dumper_179;
    nodf_module_monitor module_monitor_179;
    nodf_module_intf module_intf_180(clock,reset);
    assign module_intf_180.ap_start = 1'b0;
    assign module_intf_180.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9439.ap_ready;
    assign module_intf_180.ap_done = 1'b0;
    assign module_intf_180.ap_continue = 1'b0;
    assign module_intf_180.finish = finish;
    csv_file_dump mstatus_csv_dumper_180;
    nodf_module_monitor module_monitor_180;
    nodf_module_intf module_intf_181(clock,reset);
    assign module_intf_181.ap_start = 1'b0;
    assign module_intf_181.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9446.ap_ready;
    assign module_intf_181.ap_done = 1'b0;
    assign module_intf_181.ap_continue = 1'b0;
    assign module_intf_181.finish = finish;
    csv_file_dump mstatus_csv_dumper_181;
    nodf_module_monitor module_monitor_181;
    nodf_module_intf module_intf_182(clock,reset);
    assign module_intf_182.ap_start = 1'b0;
    assign module_intf_182.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9453.ap_ready;
    assign module_intf_182.ap_done = 1'b0;
    assign module_intf_182.ap_continue = 1'b0;
    assign module_intf_182.finish = finish;
    csv_file_dump mstatus_csv_dumper_182;
    nodf_module_monitor module_monitor_182;
    nodf_module_intf module_intf_183(clock,reset);
    assign module_intf_183.ap_start = 1'b0;
    assign module_intf_183.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9460.ap_ready;
    assign module_intf_183.ap_done = 1'b0;
    assign module_intf_183.ap_continue = 1'b0;
    assign module_intf_183.finish = finish;
    csv_file_dump mstatus_csv_dumper_183;
    nodf_module_monitor module_monitor_183;
    nodf_module_intf module_intf_184(clock,reset);
    assign module_intf_184.ap_start = 1'b0;
    assign module_intf_184.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9467.ap_ready;
    assign module_intf_184.ap_done = 1'b0;
    assign module_intf_184.ap_continue = 1'b0;
    assign module_intf_184.finish = finish;
    csv_file_dump mstatus_csv_dumper_184;
    nodf_module_monitor module_monitor_184;
    nodf_module_intf module_intf_185(clock,reset);
    assign module_intf_185.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.ap_start;
    assign module_intf_185.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.ap_ready;
    assign module_intf_185.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.ap_done;
    assign module_intf_185.ap_continue = 1'b1;
    assign module_intf_185.finish = finish;
    csv_file_dump mstatus_csv_dumper_185;
    nodf_module_monitor module_monitor_185;
    nodf_module_intf module_intf_186(clock,reset);
    assign module_intf_186.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_start;
    assign module_intf_186.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_ready;
    assign module_intf_186.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_done;
    assign module_intf_186.ap_continue = 1'b1;
    assign module_intf_186.finish = finish;
    csv_file_dump mstatus_csv_dumper_186;
    nodf_module_monitor module_monitor_186;
    nodf_module_intf module_intf_187(clock,reset);
    assign module_intf_187.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_start;
    assign module_intf_187.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_ready;
    assign module_intf_187.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_done;
    assign module_intf_187.ap_continue = 1'b1;
    assign module_intf_187.finish = finish;
    csv_file_dump mstatus_csv_dumper_187;
    nodf_module_monitor module_monitor_187;
    nodf_module_intf module_intf_188(clock,reset);
    assign module_intf_188.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_start;
    assign module_intf_188.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_ready;
    assign module_intf_188.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_done;
    assign module_intf_188.ap_continue = 1'b1;
    assign module_intf_188.finish = finish;
    csv_file_dump mstatus_csv_dumper_188;
    nodf_module_monitor module_monitor_188;
    nodf_module_intf module_intf_189(clock,reset);
    assign module_intf_189.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_start;
    assign module_intf_189.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_ready;
    assign module_intf_189.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_done;
    assign module_intf_189.ap_continue = 1'b1;
    assign module_intf_189.finish = finish;
    csv_file_dump mstatus_csv_dumper_189;
    nodf_module_monitor module_monitor_189;
    nodf_module_intf module_intf_190(clock,reset);
    assign module_intf_190.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_start;
    assign module_intf_190.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_ready;
    assign module_intf_190.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_makePatch_alignedToLine_1_fu_38373.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_done;
    assign module_intf_190.ap_continue = 1'b1;
    assign module_intf_190.finish = finish;
    csv_file_dump mstatus_csv_dumper_190;
    nodf_module_monitor module_monitor_190;
    nodf_module_intf module_intf_191(clock,reset);
    assign module_intf_191.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_delete_patch_fu_41581.ap_start;
    assign module_intf_191.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_delete_patch_fu_41581.ap_ready;
    assign module_intf_191.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_delete_patch_fu_41581.ap_done;
    assign module_intf_191.ap_continue = 1'b1;
    assign module_intf_191.finish = finish;
    csv_file_dump mstatus_csv_dumper_191;
    nodf_module_monitor module_monitor_191;
    nodf_module_intf module_intf_192(clock,reset);
    assign module_intf_192.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_delete_patch_fu_41581.grp_delete_patch_patches_parameters_fu_10118.ap_start;
    assign module_intf_192.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_delete_patch_fu_41581.grp_delete_patch_patches_parameters_fu_10118.ap_ready;
    assign module_intf_192.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_delete_patch_fu_41581.grp_delete_patch_patches_parameters_fu_10118.ap_done;
    assign module_intf_192.ap_continue = 1'b1;
    assign module_intf_192.finish = finish;
    csv_file_dump mstatus_csv_dumper_192;
    nodf_module_monitor module_monitor_192;
    nodf_module_intf module_intf_193(clock,reset);
    assign module_intf_193.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.ap_start;
    assign module_intf_193.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.ap_ready;
    assign module_intf_193.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.ap_done;
    assign module_intf_193.ap_continue = 1'b1;
    assign module_intf_193.finish = finish;
    csv_file_dump mstatus_csv_dumper_193;
    nodf_module_monitor module_monitor_193;
    nodf_module_intf module_intf_194(clock,reset);
    assign module_intf_194.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_495.ap_start;
    assign module_intf_194.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_495.ap_ready;
    assign module_intf_194.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_495.ap_done;
    assign module_intf_194.ap_continue = 1'b1;
    assign module_intf_194.finish = finish;
    csv_file_dump mstatus_csv_dumper_194;
    nodf_module_monitor module_monitor_194;
    nodf_module_intf module_intf_195(clock,reset);
    assign module_intf_195.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_509.ap_start;
    assign module_intf_195.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_509.ap_ready;
    assign module_intf_195.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_509.ap_done;
    assign module_intf_195.ap_continue = 1'b1;
    assign module_intf_195.finish = finish;
    csv_file_dump mstatus_csv_dumper_195;
    nodf_module_monitor module_monitor_195;
    nodf_module_intf module_intf_196(clock,reset);
    assign module_intf_196.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_523.ap_start;
    assign module_intf_196.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_523.ap_ready;
    assign module_intf_196.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_523.ap_done;
    assign module_intf_196.ap_continue = 1'b1;
    assign module_intf_196.finish = finish;
    csv_file_dump mstatus_csv_dumper_196;
    nodf_module_monitor module_monitor_196;
    nodf_module_intf module_intf_197(clock,reset);
    assign module_intf_197.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_537.ap_start;
    assign module_intf_197.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_537.ap_ready;
    assign module_intf_197.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_537.ap_done;
    assign module_intf_197.ap_continue = 1'b1;
    assign module_intf_197.finish = finish;
    csv_file_dump mstatus_csv_dumper_197;
    nodf_module_monitor module_monitor_197;
    nodf_module_intf module_intf_198(clock,reset);
    assign module_intf_198.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_551.ap_start;
    assign module_intf_198.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_551.ap_ready;
    assign module_intf_198.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_551.ap_done;
    assign module_intf_198.ap_continue = 1'b1;
    assign module_intf_198.finish = finish;
    csv_file_dump mstatus_csv_dumper_198;
    nodf_module_monitor module_monitor_198;
    nodf_module_intf module_intf_199(clock,reset);
    assign module_intf_199.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_565.ap_start;
    assign module_intf_199.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_565.ap_ready;
    assign module_intf_199.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_565.ap_done;
    assign module_intf_199.ap_continue = 1'b1;
    assign module_intf_199.finish = finish;
    csv_file_dump mstatus_csv_dumper_199;
    nodf_module_monitor module_monitor_199;
    nodf_module_intf module_intf_200(clock,reset);
    assign module_intf_200.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_579.ap_start;
    assign module_intf_200.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_579.ap_ready;
    assign module_intf_200.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_579.ap_done;
    assign module_intf_200.ap_continue = 1'b1;
    assign module_intf_200.finish = finish;
    csv_file_dump mstatus_csv_dumper_200;
    nodf_module_monitor module_monitor_200;
    nodf_module_intf module_intf_201(clock,reset);
    assign module_intf_201.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_593.ap_start;
    assign module_intf_201.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_593.ap_ready;
    assign module_intf_201.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_593.ap_done;
    assign module_intf_201.ap_continue = 1'b1;
    assign module_intf_201.finish = finish;
    csv_file_dump mstatus_csv_dumper_201;
    nodf_module_monitor module_monitor_201;
    nodf_module_intf module_intf_202(clock,reset);
    assign module_intf_202.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_607.ap_start;
    assign module_intf_202.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_607.ap_ready;
    assign module_intf_202.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_607.ap_done;
    assign module_intf_202.ap_continue = 1'b1;
    assign module_intf_202.finish = finish;
    csv_file_dump mstatus_csv_dumper_202;
    nodf_module_monitor module_monitor_202;
    nodf_module_intf module_intf_203(clock,reset);
    assign module_intf_203.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_621.ap_start;
    assign module_intf_203.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_621.ap_ready;
    assign module_intf_203.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_621.ap_done;
    assign module_intf_203.ap_continue = 1'b1;
    assign module_intf_203.finish = finish;
    csv_file_dump mstatus_csv_dumper_203;
    nodf_module_monitor module_monitor_203;
    nodf_module_intf module_intf_204(clock,reset);
    assign module_intf_204.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_635.ap_start;
    assign module_intf_204.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_635.ap_ready;
    assign module_intf_204.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_635.ap_done;
    assign module_intf_204.ap_continue = 1'b1;
    assign module_intf_204.finish = finish;
    csv_file_dump mstatus_csv_dumper_204;
    nodf_module_monitor module_monitor_204;
    nodf_module_intf module_intf_205(clock,reset);
    assign module_intf_205.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_649.ap_start;
    assign module_intf_205.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_649.ap_ready;
    assign module_intf_205.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_649.ap_done;
    assign module_intf_205.ap_continue = 1'b1;
    assign module_intf_205.finish = finish;
    csv_file_dump mstatus_csv_dumper_205;
    nodf_module_monitor module_monitor_205;
    nodf_module_intf module_intf_206(clock,reset);
    assign module_intf_206.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_663.ap_start;
    assign module_intf_206.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_663.ap_ready;
    assign module_intf_206.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_663.ap_done;
    assign module_intf_206.ap_continue = 1'b1;
    assign module_intf_206.finish = finish;
    csv_file_dump mstatus_csv_dumper_206;
    nodf_module_monitor module_monitor_206;
    nodf_module_intf module_intf_207(clock,reset);
    assign module_intf_207.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_677.ap_start;
    assign module_intf_207.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_677.ap_ready;
    assign module_intf_207.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_677.ap_done;
    assign module_intf_207.ap_continue = 1'b1;
    assign module_intf_207.finish = finish;
    csv_file_dump mstatus_csv_dumper_207;
    nodf_module_monitor module_monitor_207;
    nodf_module_intf module_intf_208(clock,reset);
    assign module_intf_208.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_691.ap_start;
    assign module_intf_208.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_691.ap_ready;
    assign module_intf_208.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_691.ap_done;
    assign module_intf_208.ap_continue = 1'b1;
    assign module_intf_208.finish = finish;
    csv_file_dump mstatus_csv_dumper_208;
    nodf_module_monitor module_monitor_208;
    nodf_module_intf module_intf_209(clock,reset);
    assign module_intf_209.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_705.ap_start;
    assign module_intf_209.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_705.ap_ready;
    assign module_intf_209.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makeThirdPatch_fu_39688.grp_getShadows_fu_42767.grp_straightLineProjectorFromLayerIJtoK_fu_705.ap_done;
    assign module_intf_209.ap_continue = 1'b1;
    assign module_intf_209.finish = finish;
    csv_file_dump mstatus_csv_dumper_209;
    nodf_module_monitor module_monitor_209;
    nodf_module_intf module_intf_210(clock,reset);
    assign module_intf_210.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.ap_start;
    assign module_intf_210.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.ap_ready;
    assign module_intf_210.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.ap_done;
    assign module_intf_210.ap_continue = 1'b1;
    assign module_intf_210.finish = finish;
    csv_file_dump mstatus_csv_dumper_210;
    nodf_module_monitor module_monitor_210;
    nodf_module_intf module_intf_211(clock,reset);
    assign module_intf_211.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_makeSuperPoint_alignedToLine_fu_23088.ap_start;
    assign module_intf_211.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_makeSuperPoint_alignedToLine_fu_23088.ap_ready;
    assign module_intf_211.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_makeSuperPoint_alignedToLine_fu_23088.ap_done;
    assign module_intf_211.ap_continue = 1'b1;
    assign module_intf_211.finish = finish;
    csv_file_dump mstatus_csv_dumper_211;
    nodf_module_monitor module_monitor_211;
    nodf_module_intf module_intf_212(clock,reset);
    assign module_intf_212.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_makeSuperPoint_alignedToLine_fu_23088.grp_mSP_findBounds_fu_21921.ap_start;
    assign module_intf_212.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_makeSuperPoint_alignedToLine_fu_23088.grp_mSP_findBounds_fu_21921.ap_ready;
    assign module_intf_212.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_makeSuperPoint_alignedToLine_fu_23088.grp_mSP_findBounds_fu_21921.ap_done;
    assign module_intf_212.ap_continue = 1'b1;
    assign module_intf_212.finish = finish;
    csv_file_dump mstatus_csv_dumper_212;
    nodf_module_monitor module_monitor_212;
    nodf_module_intf module_intf_213(clock,reset);
    assign module_intf_213.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.ap_start;
    assign module_intf_213.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.ap_ready;
    assign module_intf_213.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.ap_done;
    assign module_intf_213.ap_continue = 1'b1;
    assign module_intf_213.finish = finish;
    csv_file_dump mstatus_csv_dumper_213;
    nodf_module_monitor module_monitor_213;
    nodf_module_intf module_intf_214(clock,reset);
    assign module_intf_214.ap_start = 1'b0;
    assign module_intf_214.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_add_patch_patches_parameters_fu_8850.ap_ready;
    assign module_intf_214.ap_done = 1'b0;
    assign module_intf_214.ap_continue = 1'b0;
    assign module_intf_214.finish = finish;
    csv_file_dump mstatus_csv_dumper_214;
    nodf_module_monitor module_monitor_214;
    nodf_module_intf module_intf_215(clock,reset);
    assign module_intf_215.ap_start = 1'b0;
    assign module_intf_215.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8914.ap_ready;
    assign module_intf_215.ap_done = 1'b0;
    assign module_intf_215.ap_continue = 1'b0;
    assign module_intf_215.finish = finish;
    csv_file_dump mstatus_csv_dumper_215;
    nodf_module_monitor module_monitor_215;
    nodf_module_intf module_intf_216(clock,reset);
    assign module_intf_216.ap_start = 1'b0;
    assign module_intf_216.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8921.ap_ready;
    assign module_intf_216.ap_done = 1'b0;
    assign module_intf_216.ap_continue = 1'b0;
    assign module_intf_216.finish = finish;
    csv_file_dump mstatus_csv_dumper_216;
    nodf_module_monitor module_monitor_216;
    nodf_module_intf module_intf_217(clock,reset);
    assign module_intf_217.ap_start = 1'b0;
    assign module_intf_217.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8928.ap_ready;
    assign module_intf_217.ap_done = 1'b0;
    assign module_intf_217.ap_continue = 1'b0;
    assign module_intf_217.finish = finish;
    csv_file_dump mstatus_csv_dumper_217;
    nodf_module_monitor module_monitor_217;
    nodf_module_intf module_intf_218(clock,reset);
    assign module_intf_218.ap_start = 1'b0;
    assign module_intf_218.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8935.ap_ready;
    assign module_intf_218.ap_done = 1'b0;
    assign module_intf_218.ap_continue = 1'b0;
    assign module_intf_218.finish = finish;
    csv_file_dump mstatus_csv_dumper_218;
    nodf_module_monitor module_monitor_218;
    nodf_module_intf module_intf_219(clock,reset);
    assign module_intf_219.ap_start = 1'b0;
    assign module_intf_219.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8942.ap_ready;
    assign module_intf_219.ap_done = 1'b0;
    assign module_intf_219.ap_continue = 1'b0;
    assign module_intf_219.finish = finish;
    csv_file_dump mstatus_csv_dumper_219;
    nodf_module_monitor module_monitor_219;
    nodf_module_intf module_intf_220(clock,reset);
    assign module_intf_220.ap_start = 1'b0;
    assign module_intf_220.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8949.ap_ready;
    assign module_intf_220.ap_done = 1'b0;
    assign module_intf_220.ap_continue = 1'b0;
    assign module_intf_220.finish = finish;
    csv_file_dump mstatus_csv_dumper_220;
    nodf_module_monitor module_monitor_220;
    nodf_module_intf module_intf_221(clock,reset);
    assign module_intf_221.ap_start = 1'b0;
    assign module_intf_221.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8956.ap_ready;
    assign module_intf_221.ap_done = 1'b0;
    assign module_intf_221.ap_continue = 1'b0;
    assign module_intf_221.finish = finish;
    csv_file_dump mstatus_csv_dumper_221;
    nodf_module_monitor module_monitor_221;
    nodf_module_intf module_intf_222(clock,reset);
    assign module_intf_222.ap_start = 1'b0;
    assign module_intf_222.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8963.ap_ready;
    assign module_intf_222.ap_done = 1'b0;
    assign module_intf_222.ap_continue = 1'b0;
    assign module_intf_222.finish = finish;
    csv_file_dump mstatus_csv_dumper_222;
    nodf_module_monitor module_monitor_222;
    nodf_module_intf module_intf_223(clock,reset);
    assign module_intf_223.ap_start = 1'b0;
    assign module_intf_223.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8970.ap_ready;
    assign module_intf_223.ap_done = 1'b0;
    assign module_intf_223.ap_continue = 1'b0;
    assign module_intf_223.finish = finish;
    csv_file_dump mstatus_csv_dumper_223;
    nodf_module_monitor module_monitor_223;
    nodf_module_intf module_intf_224(clock,reset);
    assign module_intf_224.ap_start = 1'b0;
    assign module_intf_224.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8977.ap_ready;
    assign module_intf_224.ap_done = 1'b0;
    assign module_intf_224.ap_continue = 1'b0;
    assign module_intf_224.finish = finish;
    csv_file_dump mstatus_csv_dumper_224;
    nodf_module_monitor module_monitor_224;
    nodf_module_intf module_intf_225(clock,reset);
    assign module_intf_225.ap_start = 1'b0;
    assign module_intf_225.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8984.ap_ready;
    assign module_intf_225.ap_done = 1'b0;
    assign module_intf_225.ap_continue = 1'b0;
    assign module_intf_225.finish = finish;
    csv_file_dump mstatus_csv_dumper_225;
    nodf_module_monitor module_monitor_225;
    nodf_module_intf module_intf_226(clock,reset);
    assign module_intf_226.ap_start = 1'b0;
    assign module_intf_226.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8991.ap_ready;
    assign module_intf_226.ap_done = 1'b0;
    assign module_intf_226.ap_continue = 1'b0;
    assign module_intf_226.finish = finish;
    csv_file_dump mstatus_csv_dumper_226;
    nodf_module_monitor module_monitor_226;
    nodf_module_intf module_intf_227(clock,reset);
    assign module_intf_227.ap_start = 1'b0;
    assign module_intf_227.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_8998.ap_ready;
    assign module_intf_227.ap_done = 1'b0;
    assign module_intf_227.ap_continue = 1'b0;
    assign module_intf_227.finish = finish;
    csv_file_dump mstatus_csv_dumper_227;
    nodf_module_monitor module_monitor_227;
    nodf_module_intf module_intf_228(clock,reset);
    assign module_intf_228.ap_start = 1'b0;
    assign module_intf_228.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9005.ap_ready;
    assign module_intf_228.ap_done = 1'b0;
    assign module_intf_228.ap_continue = 1'b0;
    assign module_intf_228.finish = finish;
    csv_file_dump mstatus_csv_dumper_228;
    nodf_module_monitor module_monitor_228;
    nodf_module_intf module_intf_229(clock,reset);
    assign module_intf_229.ap_start = 1'b0;
    assign module_intf_229.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9012.ap_ready;
    assign module_intf_229.ap_done = 1'b0;
    assign module_intf_229.ap_continue = 1'b0;
    assign module_intf_229.finish = finish;
    csv_file_dump mstatus_csv_dumper_229;
    nodf_module_monitor module_monitor_229;
    nodf_module_intf module_intf_230(clock,reset);
    assign module_intf_230.ap_start = 1'b0;
    assign module_intf_230.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9019.ap_ready;
    assign module_intf_230.ap_done = 1'b0;
    assign module_intf_230.ap_continue = 1'b0;
    assign module_intf_230.finish = finish;
    csv_file_dump mstatus_csv_dumper_230;
    nodf_module_monitor module_monitor_230;
    nodf_module_intf module_intf_231(clock,reset);
    assign module_intf_231.ap_start = 1'b0;
    assign module_intf_231.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9026.ap_ready;
    assign module_intf_231.ap_done = 1'b0;
    assign module_intf_231.ap_continue = 1'b0;
    assign module_intf_231.finish = finish;
    csv_file_dump mstatus_csv_dumper_231;
    nodf_module_monitor module_monitor_231;
    nodf_module_intf module_intf_232(clock,reset);
    assign module_intf_232.ap_start = 1'b0;
    assign module_intf_232.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9033.ap_ready;
    assign module_intf_232.ap_done = 1'b0;
    assign module_intf_232.ap_continue = 1'b0;
    assign module_intf_232.finish = finish;
    csv_file_dump mstatus_csv_dumper_232;
    nodf_module_monitor module_monitor_232;
    nodf_module_intf module_intf_233(clock,reset);
    assign module_intf_233.ap_start = 1'b0;
    assign module_intf_233.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9040.ap_ready;
    assign module_intf_233.ap_done = 1'b0;
    assign module_intf_233.ap_continue = 1'b0;
    assign module_intf_233.finish = finish;
    csv_file_dump mstatus_csv_dumper_233;
    nodf_module_monitor module_monitor_233;
    nodf_module_intf module_intf_234(clock,reset);
    assign module_intf_234.ap_start = 1'b0;
    assign module_intf_234.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9047.ap_ready;
    assign module_intf_234.ap_done = 1'b0;
    assign module_intf_234.ap_continue = 1'b0;
    assign module_intf_234.finish = finish;
    csv_file_dump mstatus_csv_dumper_234;
    nodf_module_monitor module_monitor_234;
    nodf_module_intf module_intf_235(clock,reset);
    assign module_intf_235.ap_start = 1'b0;
    assign module_intf_235.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9054.ap_ready;
    assign module_intf_235.ap_done = 1'b0;
    assign module_intf_235.ap_continue = 1'b0;
    assign module_intf_235.finish = finish;
    csv_file_dump mstatus_csv_dumper_235;
    nodf_module_monitor module_monitor_235;
    nodf_module_intf module_intf_236(clock,reset);
    assign module_intf_236.ap_start = 1'b0;
    assign module_intf_236.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9061.ap_ready;
    assign module_intf_236.ap_done = 1'b0;
    assign module_intf_236.ap_continue = 1'b0;
    assign module_intf_236.finish = finish;
    csv_file_dump mstatus_csv_dumper_236;
    nodf_module_monitor module_monitor_236;
    nodf_module_intf module_intf_237(clock,reset);
    assign module_intf_237.ap_start = 1'b0;
    assign module_intf_237.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9068.ap_ready;
    assign module_intf_237.ap_done = 1'b0;
    assign module_intf_237.ap_continue = 1'b0;
    assign module_intf_237.finish = finish;
    csv_file_dump mstatus_csv_dumper_237;
    nodf_module_monitor module_monitor_237;
    nodf_module_intf module_intf_238(clock,reset);
    assign module_intf_238.ap_start = 1'b0;
    assign module_intf_238.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9075.ap_ready;
    assign module_intf_238.ap_done = 1'b0;
    assign module_intf_238.ap_continue = 1'b0;
    assign module_intf_238.finish = finish;
    csv_file_dump mstatus_csv_dumper_238;
    nodf_module_monitor module_monitor_238;
    nodf_module_intf module_intf_239(clock,reset);
    assign module_intf_239.ap_start = 1'b0;
    assign module_intf_239.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9082.ap_ready;
    assign module_intf_239.ap_done = 1'b0;
    assign module_intf_239.ap_continue = 1'b0;
    assign module_intf_239.finish = finish;
    csv_file_dump mstatus_csv_dumper_239;
    nodf_module_monitor module_monitor_239;
    nodf_module_intf module_intf_240(clock,reset);
    assign module_intf_240.ap_start = 1'b0;
    assign module_intf_240.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9089.ap_ready;
    assign module_intf_240.ap_done = 1'b0;
    assign module_intf_240.ap_continue = 1'b0;
    assign module_intf_240.finish = finish;
    csv_file_dump mstatus_csv_dumper_240;
    nodf_module_monitor module_monitor_240;
    nodf_module_intf module_intf_241(clock,reset);
    assign module_intf_241.ap_start = 1'b0;
    assign module_intf_241.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9096.ap_ready;
    assign module_intf_241.ap_done = 1'b0;
    assign module_intf_241.ap_continue = 1'b0;
    assign module_intf_241.finish = finish;
    csv_file_dump mstatus_csv_dumper_241;
    nodf_module_monitor module_monitor_241;
    nodf_module_intf module_intf_242(clock,reset);
    assign module_intf_242.ap_start = 1'b0;
    assign module_intf_242.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9103.ap_ready;
    assign module_intf_242.ap_done = 1'b0;
    assign module_intf_242.ap_continue = 1'b0;
    assign module_intf_242.finish = finish;
    csv_file_dump mstatus_csv_dumper_242;
    nodf_module_monitor module_monitor_242;
    nodf_module_intf module_intf_243(clock,reset);
    assign module_intf_243.ap_start = 1'b0;
    assign module_intf_243.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9110.ap_ready;
    assign module_intf_243.ap_done = 1'b0;
    assign module_intf_243.ap_continue = 1'b0;
    assign module_intf_243.finish = finish;
    csv_file_dump mstatus_csv_dumper_243;
    nodf_module_monitor module_monitor_243;
    nodf_module_intf module_intf_244(clock,reset);
    assign module_intf_244.ap_start = 1'b0;
    assign module_intf_244.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9117.ap_ready;
    assign module_intf_244.ap_done = 1'b0;
    assign module_intf_244.ap_continue = 1'b0;
    assign module_intf_244.finish = finish;
    csv_file_dump mstatus_csv_dumper_244;
    nodf_module_monitor module_monitor_244;
    nodf_module_intf module_intf_245(clock,reset);
    assign module_intf_245.ap_start = 1'b0;
    assign module_intf_245.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9124.ap_ready;
    assign module_intf_245.ap_done = 1'b0;
    assign module_intf_245.ap_continue = 1'b0;
    assign module_intf_245.finish = finish;
    csv_file_dump mstatus_csv_dumper_245;
    nodf_module_monitor module_monitor_245;
    nodf_module_intf module_intf_246(clock,reset);
    assign module_intf_246.ap_start = 1'b0;
    assign module_intf_246.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9131.ap_ready;
    assign module_intf_246.ap_done = 1'b0;
    assign module_intf_246.ap_continue = 1'b0;
    assign module_intf_246.finish = finish;
    csv_file_dump mstatus_csv_dumper_246;
    nodf_module_monitor module_monitor_246;
    nodf_module_intf module_intf_247(clock,reset);
    assign module_intf_247.ap_start = 1'b0;
    assign module_intf_247.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9138.ap_ready;
    assign module_intf_247.ap_done = 1'b0;
    assign module_intf_247.ap_continue = 1'b0;
    assign module_intf_247.finish = finish;
    csv_file_dump mstatus_csv_dumper_247;
    nodf_module_monitor module_monitor_247;
    nodf_module_intf module_intf_248(clock,reset);
    assign module_intf_248.ap_start = 1'b0;
    assign module_intf_248.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9145.ap_ready;
    assign module_intf_248.ap_done = 1'b0;
    assign module_intf_248.ap_continue = 1'b0;
    assign module_intf_248.finish = finish;
    csv_file_dump mstatus_csv_dumper_248;
    nodf_module_monitor module_monitor_248;
    nodf_module_intf module_intf_249(clock,reset);
    assign module_intf_249.ap_start = 1'b0;
    assign module_intf_249.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9152.ap_ready;
    assign module_intf_249.ap_done = 1'b0;
    assign module_intf_249.ap_continue = 1'b0;
    assign module_intf_249.finish = finish;
    csv_file_dump mstatus_csv_dumper_249;
    nodf_module_monitor module_monitor_249;
    nodf_module_intf module_intf_250(clock,reset);
    assign module_intf_250.ap_start = 1'b0;
    assign module_intf_250.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9159.ap_ready;
    assign module_intf_250.ap_done = 1'b0;
    assign module_intf_250.ap_continue = 1'b0;
    assign module_intf_250.finish = finish;
    csv_file_dump mstatus_csv_dumper_250;
    nodf_module_monitor module_monitor_250;
    nodf_module_intf module_intf_251(clock,reset);
    assign module_intf_251.ap_start = 1'b0;
    assign module_intf_251.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9166.ap_ready;
    assign module_intf_251.ap_done = 1'b0;
    assign module_intf_251.ap_continue = 1'b0;
    assign module_intf_251.finish = finish;
    csv_file_dump mstatus_csv_dumper_251;
    nodf_module_monitor module_monitor_251;
    nodf_module_intf module_intf_252(clock,reset);
    assign module_intf_252.ap_start = 1'b0;
    assign module_intf_252.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9173.ap_ready;
    assign module_intf_252.ap_done = 1'b0;
    assign module_intf_252.ap_continue = 1'b0;
    assign module_intf_252.finish = finish;
    csv_file_dump mstatus_csv_dumper_252;
    nodf_module_monitor module_monitor_252;
    nodf_module_intf module_intf_253(clock,reset);
    assign module_intf_253.ap_start = 1'b0;
    assign module_intf_253.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9180.ap_ready;
    assign module_intf_253.ap_done = 1'b0;
    assign module_intf_253.ap_continue = 1'b0;
    assign module_intf_253.finish = finish;
    csv_file_dump mstatus_csv_dumper_253;
    nodf_module_monitor module_monitor_253;
    nodf_module_intf module_intf_254(clock,reset);
    assign module_intf_254.ap_start = 1'b0;
    assign module_intf_254.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9187.ap_ready;
    assign module_intf_254.ap_done = 1'b0;
    assign module_intf_254.ap_continue = 1'b0;
    assign module_intf_254.finish = finish;
    csv_file_dump mstatus_csv_dumper_254;
    nodf_module_monitor module_monitor_254;
    nodf_module_intf module_intf_255(clock,reset);
    assign module_intf_255.ap_start = 1'b0;
    assign module_intf_255.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9194.ap_ready;
    assign module_intf_255.ap_done = 1'b0;
    assign module_intf_255.ap_continue = 1'b0;
    assign module_intf_255.finish = finish;
    csv_file_dump mstatus_csv_dumper_255;
    nodf_module_monitor module_monitor_255;
    nodf_module_intf module_intf_256(clock,reset);
    assign module_intf_256.ap_start = 1'b0;
    assign module_intf_256.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9201.ap_ready;
    assign module_intf_256.ap_done = 1'b0;
    assign module_intf_256.ap_continue = 1'b0;
    assign module_intf_256.finish = finish;
    csv_file_dump mstatus_csv_dumper_256;
    nodf_module_monitor module_monitor_256;
    nodf_module_intf module_intf_257(clock,reset);
    assign module_intf_257.ap_start = 1'b0;
    assign module_intf_257.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9208.ap_ready;
    assign module_intf_257.ap_done = 1'b0;
    assign module_intf_257.ap_continue = 1'b0;
    assign module_intf_257.finish = finish;
    csv_file_dump mstatus_csv_dumper_257;
    nodf_module_monitor module_monitor_257;
    nodf_module_intf module_intf_258(clock,reset);
    assign module_intf_258.ap_start = 1'b0;
    assign module_intf_258.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9215.ap_ready;
    assign module_intf_258.ap_done = 1'b0;
    assign module_intf_258.ap_continue = 1'b0;
    assign module_intf_258.finish = finish;
    csv_file_dump mstatus_csv_dumper_258;
    nodf_module_monitor module_monitor_258;
    nodf_module_intf module_intf_259(clock,reset);
    assign module_intf_259.ap_start = 1'b0;
    assign module_intf_259.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9222.ap_ready;
    assign module_intf_259.ap_done = 1'b0;
    assign module_intf_259.ap_continue = 1'b0;
    assign module_intf_259.finish = finish;
    csv_file_dump mstatus_csv_dumper_259;
    nodf_module_monitor module_monitor_259;
    nodf_module_intf module_intf_260(clock,reset);
    assign module_intf_260.ap_start = 1'b0;
    assign module_intf_260.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9229.ap_ready;
    assign module_intf_260.ap_done = 1'b0;
    assign module_intf_260.ap_continue = 1'b0;
    assign module_intf_260.finish = finish;
    csv_file_dump mstatus_csv_dumper_260;
    nodf_module_monitor module_monitor_260;
    nodf_module_intf module_intf_261(clock,reset);
    assign module_intf_261.ap_start = 1'b0;
    assign module_intf_261.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9236.ap_ready;
    assign module_intf_261.ap_done = 1'b0;
    assign module_intf_261.ap_continue = 1'b0;
    assign module_intf_261.finish = finish;
    csv_file_dump mstatus_csv_dumper_261;
    nodf_module_monitor module_monitor_261;
    nodf_module_intf module_intf_262(clock,reset);
    assign module_intf_262.ap_start = 1'b0;
    assign module_intf_262.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9243.ap_ready;
    assign module_intf_262.ap_done = 1'b0;
    assign module_intf_262.ap_continue = 1'b0;
    assign module_intf_262.finish = finish;
    csv_file_dump mstatus_csv_dumper_262;
    nodf_module_monitor module_monitor_262;
    nodf_module_intf module_intf_263(clock,reset);
    assign module_intf_263.ap_start = 1'b0;
    assign module_intf_263.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9250.ap_ready;
    assign module_intf_263.ap_done = 1'b0;
    assign module_intf_263.ap_continue = 1'b0;
    assign module_intf_263.finish = finish;
    csv_file_dump mstatus_csv_dumper_263;
    nodf_module_monitor module_monitor_263;
    nodf_module_intf module_intf_264(clock,reset);
    assign module_intf_264.ap_start = 1'b0;
    assign module_intf_264.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9257.ap_ready;
    assign module_intf_264.ap_done = 1'b0;
    assign module_intf_264.ap_continue = 1'b0;
    assign module_intf_264.finish = finish;
    csv_file_dump mstatus_csv_dumper_264;
    nodf_module_monitor module_monitor_264;
    nodf_module_intf module_intf_265(clock,reset);
    assign module_intf_265.ap_start = 1'b0;
    assign module_intf_265.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9264.ap_ready;
    assign module_intf_265.ap_done = 1'b0;
    assign module_intf_265.ap_continue = 1'b0;
    assign module_intf_265.finish = finish;
    csv_file_dump mstatus_csv_dumper_265;
    nodf_module_monitor module_monitor_265;
    nodf_module_intf module_intf_266(clock,reset);
    assign module_intf_266.ap_start = 1'b0;
    assign module_intf_266.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9271.ap_ready;
    assign module_intf_266.ap_done = 1'b0;
    assign module_intf_266.ap_continue = 1'b0;
    assign module_intf_266.finish = finish;
    csv_file_dump mstatus_csv_dumper_266;
    nodf_module_monitor module_monitor_266;
    nodf_module_intf module_intf_267(clock,reset);
    assign module_intf_267.ap_start = 1'b0;
    assign module_intf_267.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9278.ap_ready;
    assign module_intf_267.ap_done = 1'b0;
    assign module_intf_267.ap_continue = 1'b0;
    assign module_intf_267.finish = finish;
    csv_file_dump mstatus_csv_dumper_267;
    nodf_module_monitor module_monitor_267;
    nodf_module_intf module_intf_268(clock,reset);
    assign module_intf_268.ap_start = 1'b0;
    assign module_intf_268.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9285.ap_ready;
    assign module_intf_268.ap_done = 1'b0;
    assign module_intf_268.ap_continue = 1'b0;
    assign module_intf_268.finish = finish;
    csv_file_dump mstatus_csv_dumper_268;
    nodf_module_monitor module_monitor_268;
    nodf_module_intf module_intf_269(clock,reset);
    assign module_intf_269.ap_start = 1'b0;
    assign module_intf_269.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9292.ap_ready;
    assign module_intf_269.ap_done = 1'b0;
    assign module_intf_269.ap_continue = 1'b0;
    assign module_intf_269.finish = finish;
    csv_file_dump mstatus_csv_dumper_269;
    nodf_module_monitor module_monitor_269;
    nodf_module_intf module_intf_270(clock,reset);
    assign module_intf_270.ap_start = 1'b0;
    assign module_intf_270.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9299.ap_ready;
    assign module_intf_270.ap_done = 1'b0;
    assign module_intf_270.ap_continue = 1'b0;
    assign module_intf_270.finish = finish;
    csv_file_dump mstatus_csv_dumper_270;
    nodf_module_monitor module_monitor_270;
    nodf_module_intf module_intf_271(clock,reset);
    assign module_intf_271.ap_start = 1'b0;
    assign module_intf_271.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9306.ap_ready;
    assign module_intf_271.ap_done = 1'b0;
    assign module_intf_271.ap_continue = 1'b0;
    assign module_intf_271.finish = finish;
    csv_file_dump mstatus_csv_dumper_271;
    nodf_module_monitor module_monitor_271;
    nodf_module_intf module_intf_272(clock,reset);
    assign module_intf_272.ap_start = 1'b0;
    assign module_intf_272.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9313.ap_ready;
    assign module_intf_272.ap_done = 1'b0;
    assign module_intf_272.ap_continue = 1'b0;
    assign module_intf_272.finish = finish;
    csv_file_dump mstatus_csv_dumper_272;
    nodf_module_monitor module_monitor_272;
    nodf_module_intf module_intf_273(clock,reset);
    assign module_intf_273.ap_start = 1'b0;
    assign module_intf_273.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9320.ap_ready;
    assign module_intf_273.ap_done = 1'b0;
    assign module_intf_273.ap_continue = 1'b0;
    assign module_intf_273.finish = finish;
    csv_file_dump mstatus_csv_dumper_273;
    nodf_module_monitor module_monitor_273;
    nodf_module_intf module_intf_274(clock,reset);
    assign module_intf_274.ap_start = 1'b0;
    assign module_intf_274.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9327.ap_ready;
    assign module_intf_274.ap_done = 1'b0;
    assign module_intf_274.ap_continue = 1'b0;
    assign module_intf_274.finish = finish;
    csv_file_dump mstatus_csv_dumper_274;
    nodf_module_monitor module_monitor_274;
    nodf_module_intf module_intf_275(clock,reset);
    assign module_intf_275.ap_start = 1'b0;
    assign module_intf_275.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9334.ap_ready;
    assign module_intf_275.ap_done = 1'b0;
    assign module_intf_275.ap_continue = 1'b0;
    assign module_intf_275.finish = finish;
    csv_file_dump mstatus_csv_dumper_275;
    nodf_module_monitor module_monitor_275;
    nodf_module_intf module_intf_276(clock,reset);
    assign module_intf_276.ap_start = 1'b0;
    assign module_intf_276.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9341.ap_ready;
    assign module_intf_276.ap_done = 1'b0;
    assign module_intf_276.ap_continue = 1'b0;
    assign module_intf_276.finish = finish;
    csv_file_dump mstatus_csv_dumper_276;
    nodf_module_monitor module_monitor_276;
    nodf_module_intf module_intf_277(clock,reset);
    assign module_intf_277.ap_start = 1'b0;
    assign module_intf_277.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9348.ap_ready;
    assign module_intf_277.ap_done = 1'b0;
    assign module_intf_277.ap_continue = 1'b0;
    assign module_intf_277.finish = finish;
    csv_file_dump mstatus_csv_dumper_277;
    nodf_module_monitor module_monitor_277;
    nodf_module_intf module_intf_278(clock,reset);
    assign module_intf_278.ap_start = 1'b0;
    assign module_intf_278.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9355.ap_ready;
    assign module_intf_278.ap_done = 1'b0;
    assign module_intf_278.ap_continue = 1'b0;
    assign module_intf_278.finish = finish;
    csv_file_dump mstatus_csv_dumper_278;
    nodf_module_monitor module_monitor_278;
    nodf_module_intf module_intf_279(clock,reset);
    assign module_intf_279.ap_start = 1'b0;
    assign module_intf_279.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9362.ap_ready;
    assign module_intf_279.ap_done = 1'b0;
    assign module_intf_279.ap_continue = 1'b0;
    assign module_intf_279.finish = finish;
    csv_file_dump mstatus_csv_dumper_279;
    nodf_module_monitor module_monitor_279;
    nodf_module_intf module_intf_280(clock,reset);
    assign module_intf_280.ap_start = 1'b0;
    assign module_intf_280.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9369.ap_ready;
    assign module_intf_280.ap_done = 1'b0;
    assign module_intf_280.ap_continue = 1'b0;
    assign module_intf_280.finish = finish;
    csv_file_dump mstatus_csv_dumper_280;
    nodf_module_monitor module_monitor_280;
    nodf_module_intf module_intf_281(clock,reset);
    assign module_intf_281.ap_start = 1'b0;
    assign module_intf_281.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9376.ap_ready;
    assign module_intf_281.ap_done = 1'b0;
    assign module_intf_281.ap_continue = 1'b0;
    assign module_intf_281.finish = finish;
    csv_file_dump mstatus_csv_dumper_281;
    nodf_module_monitor module_monitor_281;
    nodf_module_intf module_intf_282(clock,reset);
    assign module_intf_282.ap_start = 1'b0;
    assign module_intf_282.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9383.ap_ready;
    assign module_intf_282.ap_done = 1'b0;
    assign module_intf_282.ap_continue = 1'b0;
    assign module_intf_282.finish = finish;
    csv_file_dump mstatus_csv_dumper_282;
    nodf_module_monitor module_monitor_282;
    nodf_module_intf module_intf_283(clock,reset);
    assign module_intf_283.ap_start = 1'b0;
    assign module_intf_283.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9390.ap_ready;
    assign module_intf_283.ap_done = 1'b0;
    assign module_intf_283.ap_continue = 1'b0;
    assign module_intf_283.finish = finish;
    csv_file_dump mstatus_csv_dumper_283;
    nodf_module_monitor module_monitor_283;
    nodf_module_intf module_intf_284(clock,reset);
    assign module_intf_284.ap_start = 1'b0;
    assign module_intf_284.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9397.ap_ready;
    assign module_intf_284.ap_done = 1'b0;
    assign module_intf_284.ap_continue = 1'b0;
    assign module_intf_284.finish = finish;
    csv_file_dump mstatus_csv_dumper_284;
    nodf_module_monitor module_monitor_284;
    nodf_module_intf module_intf_285(clock,reset);
    assign module_intf_285.ap_start = 1'b0;
    assign module_intf_285.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9404.ap_ready;
    assign module_intf_285.ap_done = 1'b0;
    assign module_intf_285.ap_continue = 1'b0;
    assign module_intf_285.finish = finish;
    csv_file_dump mstatus_csv_dumper_285;
    nodf_module_monitor module_monitor_285;
    nodf_module_intf module_intf_286(clock,reset);
    assign module_intf_286.ap_start = 1'b0;
    assign module_intf_286.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9411.ap_ready;
    assign module_intf_286.ap_done = 1'b0;
    assign module_intf_286.ap_continue = 1'b0;
    assign module_intf_286.finish = finish;
    csv_file_dump mstatus_csv_dumper_286;
    nodf_module_monitor module_monitor_286;
    nodf_module_intf module_intf_287(clock,reset);
    assign module_intf_287.ap_start = 1'b0;
    assign module_intf_287.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9418.ap_ready;
    assign module_intf_287.ap_done = 1'b0;
    assign module_intf_287.ap_continue = 1'b0;
    assign module_intf_287.finish = finish;
    csv_file_dump mstatus_csv_dumper_287;
    nodf_module_monitor module_monitor_287;
    nodf_module_intf module_intf_288(clock,reset);
    assign module_intf_288.ap_start = 1'b0;
    assign module_intf_288.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9425.ap_ready;
    assign module_intf_288.ap_done = 1'b0;
    assign module_intf_288.ap_continue = 1'b0;
    assign module_intf_288.finish = finish;
    csv_file_dump mstatus_csv_dumper_288;
    nodf_module_monitor module_monitor_288;
    nodf_module_intf module_intf_289(clock,reset);
    assign module_intf_289.ap_start = 1'b0;
    assign module_intf_289.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9432.ap_ready;
    assign module_intf_289.ap_done = 1'b0;
    assign module_intf_289.ap_continue = 1'b0;
    assign module_intf_289.finish = finish;
    csv_file_dump mstatus_csv_dumper_289;
    nodf_module_monitor module_monitor_289;
    nodf_module_intf module_intf_290(clock,reset);
    assign module_intf_290.ap_start = 1'b0;
    assign module_intf_290.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9439.ap_ready;
    assign module_intf_290.ap_done = 1'b0;
    assign module_intf_290.ap_continue = 1'b0;
    assign module_intf_290.finish = finish;
    csv_file_dump mstatus_csv_dumper_290;
    nodf_module_monitor module_monitor_290;
    nodf_module_intf module_intf_291(clock,reset);
    assign module_intf_291.ap_start = 1'b0;
    assign module_intf_291.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9446.ap_ready;
    assign module_intf_291.ap_done = 1'b0;
    assign module_intf_291.ap_continue = 1'b0;
    assign module_intf_291.finish = finish;
    csv_file_dump mstatus_csv_dumper_291;
    nodf_module_monitor module_monitor_291;
    nodf_module_intf module_intf_292(clock,reset);
    assign module_intf_292.ap_start = 1'b0;
    assign module_intf_292.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9453.ap_ready;
    assign module_intf_292.ap_done = 1'b0;
    assign module_intf_292.ap_continue = 1'b0;
    assign module_intf_292.finish = finish;
    csv_file_dump mstatus_csv_dumper_292;
    nodf_module_monitor module_monitor_292;
    nodf_module_intf module_intf_293(clock,reset);
    assign module_intf_293.ap_start = 1'b0;
    assign module_intf_293.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9460.ap_ready;
    assign module_intf_293.ap_done = 1'b0;
    assign module_intf_293.ap_continue = 1'b0;
    assign module_intf_293.finish = finish;
    csv_file_dump mstatus_csv_dumper_293;
    nodf_module_monitor module_monitor_293;
    nodf_module_intf module_intf_294(clock,reset);
    assign module_intf_294.ap_start = 1'b0;
    assign module_intf_294.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_fu_42900.grp_add_patch_fu_28558.grp_encodeCoordinates_fu_9467.ap_ready;
    assign module_intf_294.ap_done = 1'b0;
    assign module_intf_294.ap_continue = 1'b0;
    assign module_intf_294.finish = finish;
    csv_file_dump mstatus_csv_dumper_294;
    nodf_module_monitor module_monitor_294;
    nodf_module_intf module_intf_295(clock,reset);
    assign module_intf_295.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.ap_start;
    assign module_intf_295.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.ap_ready;
    assign module_intf_295.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.ap_done;
    assign module_intf_295.ap_continue = 1'b1;
    assign module_intf_295.finish = finish;
    csv_file_dump mstatus_csv_dumper_295;
    nodf_module_monitor module_monitor_295;
    nodf_module_intf module_intf_296(clock,reset);
    assign module_intf_296.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_makeSuperPoint_alignedToLine_1_fu_23098.ap_start;
    assign module_intf_296.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_makeSuperPoint_alignedToLine_1_fu_23098.ap_ready;
    assign module_intf_296.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_makeSuperPoint_alignedToLine_1_fu_23098.ap_done;
    assign module_intf_296.ap_continue = 1'b1;
    assign module_intf_296.finish = finish;
    csv_file_dump mstatus_csv_dumper_296;
    nodf_module_monitor module_monitor_296;
    nodf_module_intf module_intf_297(clock,reset);
    assign module_intf_297.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_makeSuperPoint_alignedToLine_1_fu_23098.grp_mSP_findBounds_fu_21935.ap_start;
    assign module_intf_297.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_makeSuperPoint_alignedToLine_1_fu_23098.grp_mSP_findBounds_fu_21935.ap_ready;
    assign module_intf_297.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_makeSuperPoint_alignedToLine_1_fu_23098.grp_mSP_findBounds_fu_21935.ap_done;
    assign module_intf_297.ap_continue = 1'b1;
    assign module_intf_297.finish = finish;
    csv_file_dump mstatus_csv_dumper_297;
    nodf_module_monitor module_monitor_297;
    nodf_module_intf module_intf_298(clock,reset);
    assign module_intf_298.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.ap_start;
    assign module_intf_298.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.ap_ready;
    assign module_intf_298.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.ap_done;
    assign module_intf_298.ap_continue = 1'b1;
    assign module_intf_298.finish = finish;
    csv_file_dump mstatus_csv_dumper_298;
    nodf_module_monitor module_monitor_298;
    nodf_module_intf module_intf_299(clock,reset);
    assign module_intf_299.ap_start = 1'b0;
    assign module_intf_299.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_add_patch_patches_parameters_fu_8850.ap_ready;
    assign module_intf_299.ap_done = 1'b0;
    assign module_intf_299.ap_continue = 1'b0;
    assign module_intf_299.finish = finish;
    csv_file_dump mstatus_csv_dumper_299;
    nodf_module_monitor module_monitor_299;
    nodf_module_intf module_intf_300(clock,reset);
    assign module_intf_300.ap_start = 1'b0;
    assign module_intf_300.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8914.ap_ready;
    assign module_intf_300.ap_done = 1'b0;
    assign module_intf_300.ap_continue = 1'b0;
    assign module_intf_300.finish = finish;
    csv_file_dump mstatus_csv_dumper_300;
    nodf_module_monitor module_monitor_300;
    nodf_module_intf module_intf_301(clock,reset);
    assign module_intf_301.ap_start = 1'b0;
    assign module_intf_301.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8921.ap_ready;
    assign module_intf_301.ap_done = 1'b0;
    assign module_intf_301.ap_continue = 1'b0;
    assign module_intf_301.finish = finish;
    csv_file_dump mstatus_csv_dumper_301;
    nodf_module_monitor module_monitor_301;
    nodf_module_intf module_intf_302(clock,reset);
    assign module_intf_302.ap_start = 1'b0;
    assign module_intf_302.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8928.ap_ready;
    assign module_intf_302.ap_done = 1'b0;
    assign module_intf_302.ap_continue = 1'b0;
    assign module_intf_302.finish = finish;
    csv_file_dump mstatus_csv_dumper_302;
    nodf_module_monitor module_monitor_302;
    nodf_module_intf module_intf_303(clock,reset);
    assign module_intf_303.ap_start = 1'b0;
    assign module_intf_303.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8935.ap_ready;
    assign module_intf_303.ap_done = 1'b0;
    assign module_intf_303.ap_continue = 1'b0;
    assign module_intf_303.finish = finish;
    csv_file_dump mstatus_csv_dumper_303;
    nodf_module_monitor module_monitor_303;
    nodf_module_intf module_intf_304(clock,reset);
    assign module_intf_304.ap_start = 1'b0;
    assign module_intf_304.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8942.ap_ready;
    assign module_intf_304.ap_done = 1'b0;
    assign module_intf_304.ap_continue = 1'b0;
    assign module_intf_304.finish = finish;
    csv_file_dump mstatus_csv_dumper_304;
    nodf_module_monitor module_monitor_304;
    nodf_module_intf module_intf_305(clock,reset);
    assign module_intf_305.ap_start = 1'b0;
    assign module_intf_305.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8949.ap_ready;
    assign module_intf_305.ap_done = 1'b0;
    assign module_intf_305.ap_continue = 1'b0;
    assign module_intf_305.finish = finish;
    csv_file_dump mstatus_csv_dumper_305;
    nodf_module_monitor module_monitor_305;
    nodf_module_intf module_intf_306(clock,reset);
    assign module_intf_306.ap_start = 1'b0;
    assign module_intf_306.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8956.ap_ready;
    assign module_intf_306.ap_done = 1'b0;
    assign module_intf_306.ap_continue = 1'b0;
    assign module_intf_306.finish = finish;
    csv_file_dump mstatus_csv_dumper_306;
    nodf_module_monitor module_monitor_306;
    nodf_module_intf module_intf_307(clock,reset);
    assign module_intf_307.ap_start = 1'b0;
    assign module_intf_307.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8963.ap_ready;
    assign module_intf_307.ap_done = 1'b0;
    assign module_intf_307.ap_continue = 1'b0;
    assign module_intf_307.finish = finish;
    csv_file_dump mstatus_csv_dumper_307;
    nodf_module_monitor module_monitor_307;
    nodf_module_intf module_intf_308(clock,reset);
    assign module_intf_308.ap_start = 1'b0;
    assign module_intf_308.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8970.ap_ready;
    assign module_intf_308.ap_done = 1'b0;
    assign module_intf_308.ap_continue = 1'b0;
    assign module_intf_308.finish = finish;
    csv_file_dump mstatus_csv_dumper_308;
    nodf_module_monitor module_monitor_308;
    nodf_module_intf module_intf_309(clock,reset);
    assign module_intf_309.ap_start = 1'b0;
    assign module_intf_309.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8977.ap_ready;
    assign module_intf_309.ap_done = 1'b0;
    assign module_intf_309.ap_continue = 1'b0;
    assign module_intf_309.finish = finish;
    csv_file_dump mstatus_csv_dumper_309;
    nodf_module_monitor module_monitor_309;
    nodf_module_intf module_intf_310(clock,reset);
    assign module_intf_310.ap_start = 1'b0;
    assign module_intf_310.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8984.ap_ready;
    assign module_intf_310.ap_done = 1'b0;
    assign module_intf_310.ap_continue = 1'b0;
    assign module_intf_310.finish = finish;
    csv_file_dump mstatus_csv_dumper_310;
    nodf_module_monitor module_monitor_310;
    nodf_module_intf module_intf_311(clock,reset);
    assign module_intf_311.ap_start = 1'b0;
    assign module_intf_311.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8991.ap_ready;
    assign module_intf_311.ap_done = 1'b0;
    assign module_intf_311.ap_continue = 1'b0;
    assign module_intf_311.finish = finish;
    csv_file_dump mstatus_csv_dumper_311;
    nodf_module_monitor module_monitor_311;
    nodf_module_intf module_intf_312(clock,reset);
    assign module_intf_312.ap_start = 1'b0;
    assign module_intf_312.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_8998.ap_ready;
    assign module_intf_312.ap_done = 1'b0;
    assign module_intf_312.ap_continue = 1'b0;
    assign module_intf_312.finish = finish;
    csv_file_dump mstatus_csv_dumper_312;
    nodf_module_monitor module_monitor_312;
    nodf_module_intf module_intf_313(clock,reset);
    assign module_intf_313.ap_start = 1'b0;
    assign module_intf_313.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9005.ap_ready;
    assign module_intf_313.ap_done = 1'b0;
    assign module_intf_313.ap_continue = 1'b0;
    assign module_intf_313.finish = finish;
    csv_file_dump mstatus_csv_dumper_313;
    nodf_module_monitor module_monitor_313;
    nodf_module_intf module_intf_314(clock,reset);
    assign module_intf_314.ap_start = 1'b0;
    assign module_intf_314.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9012.ap_ready;
    assign module_intf_314.ap_done = 1'b0;
    assign module_intf_314.ap_continue = 1'b0;
    assign module_intf_314.finish = finish;
    csv_file_dump mstatus_csv_dumper_314;
    nodf_module_monitor module_monitor_314;
    nodf_module_intf module_intf_315(clock,reset);
    assign module_intf_315.ap_start = 1'b0;
    assign module_intf_315.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9019.ap_ready;
    assign module_intf_315.ap_done = 1'b0;
    assign module_intf_315.ap_continue = 1'b0;
    assign module_intf_315.finish = finish;
    csv_file_dump mstatus_csv_dumper_315;
    nodf_module_monitor module_monitor_315;
    nodf_module_intf module_intf_316(clock,reset);
    assign module_intf_316.ap_start = 1'b0;
    assign module_intf_316.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9026.ap_ready;
    assign module_intf_316.ap_done = 1'b0;
    assign module_intf_316.ap_continue = 1'b0;
    assign module_intf_316.finish = finish;
    csv_file_dump mstatus_csv_dumper_316;
    nodf_module_monitor module_monitor_316;
    nodf_module_intf module_intf_317(clock,reset);
    assign module_intf_317.ap_start = 1'b0;
    assign module_intf_317.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9033.ap_ready;
    assign module_intf_317.ap_done = 1'b0;
    assign module_intf_317.ap_continue = 1'b0;
    assign module_intf_317.finish = finish;
    csv_file_dump mstatus_csv_dumper_317;
    nodf_module_monitor module_monitor_317;
    nodf_module_intf module_intf_318(clock,reset);
    assign module_intf_318.ap_start = 1'b0;
    assign module_intf_318.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9040.ap_ready;
    assign module_intf_318.ap_done = 1'b0;
    assign module_intf_318.ap_continue = 1'b0;
    assign module_intf_318.finish = finish;
    csv_file_dump mstatus_csv_dumper_318;
    nodf_module_monitor module_monitor_318;
    nodf_module_intf module_intf_319(clock,reset);
    assign module_intf_319.ap_start = 1'b0;
    assign module_intf_319.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9047.ap_ready;
    assign module_intf_319.ap_done = 1'b0;
    assign module_intf_319.ap_continue = 1'b0;
    assign module_intf_319.finish = finish;
    csv_file_dump mstatus_csv_dumper_319;
    nodf_module_monitor module_monitor_319;
    nodf_module_intf module_intf_320(clock,reset);
    assign module_intf_320.ap_start = 1'b0;
    assign module_intf_320.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9054.ap_ready;
    assign module_intf_320.ap_done = 1'b0;
    assign module_intf_320.ap_continue = 1'b0;
    assign module_intf_320.finish = finish;
    csv_file_dump mstatus_csv_dumper_320;
    nodf_module_monitor module_monitor_320;
    nodf_module_intf module_intf_321(clock,reset);
    assign module_intf_321.ap_start = 1'b0;
    assign module_intf_321.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9061.ap_ready;
    assign module_intf_321.ap_done = 1'b0;
    assign module_intf_321.ap_continue = 1'b0;
    assign module_intf_321.finish = finish;
    csv_file_dump mstatus_csv_dumper_321;
    nodf_module_monitor module_monitor_321;
    nodf_module_intf module_intf_322(clock,reset);
    assign module_intf_322.ap_start = 1'b0;
    assign module_intf_322.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9068.ap_ready;
    assign module_intf_322.ap_done = 1'b0;
    assign module_intf_322.ap_continue = 1'b0;
    assign module_intf_322.finish = finish;
    csv_file_dump mstatus_csv_dumper_322;
    nodf_module_monitor module_monitor_322;
    nodf_module_intf module_intf_323(clock,reset);
    assign module_intf_323.ap_start = 1'b0;
    assign module_intf_323.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9075.ap_ready;
    assign module_intf_323.ap_done = 1'b0;
    assign module_intf_323.ap_continue = 1'b0;
    assign module_intf_323.finish = finish;
    csv_file_dump mstatus_csv_dumper_323;
    nodf_module_monitor module_monitor_323;
    nodf_module_intf module_intf_324(clock,reset);
    assign module_intf_324.ap_start = 1'b0;
    assign module_intf_324.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9082.ap_ready;
    assign module_intf_324.ap_done = 1'b0;
    assign module_intf_324.ap_continue = 1'b0;
    assign module_intf_324.finish = finish;
    csv_file_dump mstatus_csv_dumper_324;
    nodf_module_monitor module_monitor_324;
    nodf_module_intf module_intf_325(clock,reset);
    assign module_intf_325.ap_start = 1'b0;
    assign module_intf_325.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9089.ap_ready;
    assign module_intf_325.ap_done = 1'b0;
    assign module_intf_325.ap_continue = 1'b0;
    assign module_intf_325.finish = finish;
    csv_file_dump mstatus_csv_dumper_325;
    nodf_module_monitor module_monitor_325;
    nodf_module_intf module_intf_326(clock,reset);
    assign module_intf_326.ap_start = 1'b0;
    assign module_intf_326.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9096.ap_ready;
    assign module_intf_326.ap_done = 1'b0;
    assign module_intf_326.ap_continue = 1'b0;
    assign module_intf_326.finish = finish;
    csv_file_dump mstatus_csv_dumper_326;
    nodf_module_monitor module_monitor_326;
    nodf_module_intf module_intf_327(clock,reset);
    assign module_intf_327.ap_start = 1'b0;
    assign module_intf_327.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9103.ap_ready;
    assign module_intf_327.ap_done = 1'b0;
    assign module_intf_327.ap_continue = 1'b0;
    assign module_intf_327.finish = finish;
    csv_file_dump mstatus_csv_dumper_327;
    nodf_module_monitor module_monitor_327;
    nodf_module_intf module_intf_328(clock,reset);
    assign module_intf_328.ap_start = 1'b0;
    assign module_intf_328.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9110.ap_ready;
    assign module_intf_328.ap_done = 1'b0;
    assign module_intf_328.ap_continue = 1'b0;
    assign module_intf_328.finish = finish;
    csv_file_dump mstatus_csv_dumper_328;
    nodf_module_monitor module_monitor_328;
    nodf_module_intf module_intf_329(clock,reset);
    assign module_intf_329.ap_start = 1'b0;
    assign module_intf_329.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9117.ap_ready;
    assign module_intf_329.ap_done = 1'b0;
    assign module_intf_329.ap_continue = 1'b0;
    assign module_intf_329.finish = finish;
    csv_file_dump mstatus_csv_dumper_329;
    nodf_module_monitor module_monitor_329;
    nodf_module_intf module_intf_330(clock,reset);
    assign module_intf_330.ap_start = 1'b0;
    assign module_intf_330.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9124.ap_ready;
    assign module_intf_330.ap_done = 1'b0;
    assign module_intf_330.ap_continue = 1'b0;
    assign module_intf_330.finish = finish;
    csv_file_dump mstatus_csv_dumper_330;
    nodf_module_monitor module_monitor_330;
    nodf_module_intf module_intf_331(clock,reset);
    assign module_intf_331.ap_start = 1'b0;
    assign module_intf_331.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9131.ap_ready;
    assign module_intf_331.ap_done = 1'b0;
    assign module_intf_331.ap_continue = 1'b0;
    assign module_intf_331.finish = finish;
    csv_file_dump mstatus_csv_dumper_331;
    nodf_module_monitor module_monitor_331;
    nodf_module_intf module_intf_332(clock,reset);
    assign module_intf_332.ap_start = 1'b0;
    assign module_intf_332.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9138.ap_ready;
    assign module_intf_332.ap_done = 1'b0;
    assign module_intf_332.ap_continue = 1'b0;
    assign module_intf_332.finish = finish;
    csv_file_dump mstatus_csv_dumper_332;
    nodf_module_monitor module_monitor_332;
    nodf_module_intf module_intf_333(clock,reset);
    assign module_intf_333.ap_start = 1'b0;
    assign module_intf_333.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9145.ap_ready;
    assign module_intf_333.ap_done = 1'b0;
    assign module_intf_333.ap_continue = 1'b0;
    assign module_intf_333.finish = finish;
    csv_file_dump mstatus_csv_dumper_333;
    nodf_module_monitor module_monitor_333;
    nodf_module_intf module_intf_334(clock,reset);
    assign module_intf_334.ap_start = 1'b0;
    assign module_intf_334.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9152.ap_ready;
    assign module_intf_334.ap_done = 1'b0;
    assign module_intf_334.ap_continue = 1'b0;
    assign module_intf_334.finish = finish;
    csv_file_dump mstatus_csv_dumper_334;
    nodf_module_monitor module_monitor_334;
    nodf_module_intf module_intf_335(clock,reset);
    assign module_intf_335.ap_start = 1'b0;
    assign module_intf_335.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9159.ap_ready;
    assign module_intf_335.ap_done = 1'b0;
    assign module_intf_335.ap_continue = 1'b0;
    assign module_intf_335.finish = finish;
    csv_file_dump mstatus_csv_dumper_335;
    nodf_module_monitor module_monitor_335;
    nodf_module_intf module_intf_336(clock,reset);
    assign module_intf_336.ap_start = 1'b0;
    assign module_intf_336.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9166.ap_ready;
    assign module_intf_336.ap_done = 1'b0;
    assign module_intf_336.ap_continue = 1'b0;
    assign module_intf_336.finish = finish;
    csv_file_dump mstatus_csv_dumper_336;
    nodf_module_monitor module_monitor_336;
    nodf_module_intf module_intf_337(clock,reset);
    assign module_intf_337.ap_start = 1'b0;
    assign module_intf_337.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9173.ap_ready;
    assign module_intf_337.ap_done = 1'b0;
    assign module_intf_337.ap_continue = 1'b0;
    assign module_intf_337.finish = finish;
    csv_file_dump mstatus_csv_dumper_337;
    nodf_module_monitor module_monitor_337;
    nodf_module_intf module_intf_338(clock,reset);
    assign module_intf_338.ap_start = 1'b0;
    assign module_intf_338.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9180.ap_ready;
    assign module_intf_338.ap_done = 1'b0;
    assign module_intf_338.ap_continue = 1'b0;
    assign module_intf_338.finish = finish;
    csv_file_dump mstatus_csv_dumper_338;
    nodf_module_monitor module_monitor_338;
    nodf_module_intf module_intf_339(clock,reset);
    assign module_intf_339.ap_start = 1'b0;
    assign module_intf_339.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9187.ap_ready;
    assign module_intf_339.ap_done = 1'b0;
    assign module_intf_339.ap_continue = 1'b0;
    assign module_intf_339.finish = finish;
    csv_file_dump mstatus_csv_dumper_339;
    nodf_module_monitor module_monitor_339;
    nodf_module_intf module_intf_340(clock,reset);
    assign module_intf_340.ap_start = 1'b0;
    assign module_intf_340.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9194.ap_ready;
    assign module_intf_340.ap_done = 1'b0;
    assign module_intf_340.ap_continue = 1'b0;
    assign module_intf_340.finish = finish;
    csv_file_dump mstatus_csv_dumper_340;
    nodf_module_monitor module_monitor_340;
    nodf_module_intf module_intf_341(clock,reset);
    assign module_intf_341.ap_start = 1'b0;
    assign module_intf_341.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9201.ap_ready;
    assign module_intf_341.ap_done = 1'b0;
    assign module_intf_341.ap_continue = 1'b0;
    assign module_intf_341.finish = finish;
    csv_file_dump mstatus_csv_dumper_341;
    nodf_module_monitor module_monitor_341;
    nodf_module_intf module_intf_342(clock,reset);
    assign module_intf_342.ap_start = 1'b0;
    assign module_intf_342.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9208.ap_ready;
    assign module_intf_342.ap_done = 1'b0;
    assign module_intf_342.ap_continue = 1'b0;
    assign module_intf_342.finish = finish;
    csv_file_dump mstatus_csv_dumper_342;
    nodf_module_monitor module_monitor_342;
    nodf_module_intf module_intf_343(clock,reset);
    assign module_intf_343.ap_start = 1'b0;
    assign module_intf_343.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9215.ap_ready;
    assign module_intf_343.ap_done = 1'b0;
    assign module_intf_343.ap_continue = 1'b0;
    assign module_intf_343.finish = finish;
    csv_file_dump mstatus_csv_dumper_343;
    nodf_module_monitor module_monitor_343;
    nodf_module_intf module_intf_344(clock,reset);
    assign module_intf_344.ap_start = 1'b0;
    assign module_intf_344.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9222.ap_ready;
    assign module_intf_344.ap_done = 1'b0;
    assign module_intf_344.ap_continue = 1'b0;
    assign module_intf_344.finish = finish;
    csv_file_dump mstatus_csv_dumper_344;
    nodf_module_monitor module_monitor_344;
    nodf_module_intf module_intf_345(clock,reset);
    assign module_intf_345.ap_start = 1'b0;
    assign module_intf_345.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9229.ap_ready;
    assign module_intf_345.ap_done = 1'b0;
    assign module_intf_345.ap_continue = 1'b0;
    assign module_intf_345.finish = finish;
    csv_file_dump mstatus_csv_dumper_345;
    nodf_module_monitor module_monitor_345;
    nodf_module_intf module_intf_346(clock,reset);
    assign module_intf_346.ap_start = 1'b0;
    assign module_intf_346.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9236.ap_ready;
    assign module_intf_346.ap_done = 1'b0;
    assign module_intf_346.ap_continue = 1'b0;
    assign module_intf_346.finish = finish;
    csv_file_dump mstatus_csv_dumper_346;
    nodf_module_monitor module_monitor_346;
    nodf_module_intf module_intf_347(clock,reset);
    assign module_intf_347.ap_start = 1'b0;
    assign module_intf_347.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9243.ap_ready;
    assign module_intf_347.ap_done = 1'b0;
    assign module_intf_347.ap_continue = 1'b0;
    assign module_intf_347.finish = finish;
    csv_file_dump mstatus_csv_dumper_347;
    nodf_module_monitor module_monitor_347;
    nodf_module_intf module_intf_348(clock,reset);
    assign module_intf_348.ap_start = 1'b0;
    assign module_intf_348.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9250.ap_ready;
    assign module_intf_348.ap_done = 1'b0;
    assign module_intf_348.ap_continue = 1'b0;
    assign module_intf_348.finish = finish;
    csv_file_dump mstatus_csv_dumper_348;
    nodf_module_monitor module_monitor_348;
    nodf_module_intf module_intf_349(clock,reset);
    assign module_intf_349.ap_start = 1'b0;
    assign module_intf_349.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9257.ap_ready;
    assign module_intf_349.ap_done = 1'b0;
    assign module_intf_349.ap_continue = 1'b0;
    assign module_intf_349.finish = finish;
    csv_file_dump mstatus_csv_dumper_349;
    nodf_module_monitor module_monitor_349;
    nodf_module_intf module_intf_350(clock,reset);
    assign module_intf_350.ap_start = 1'b0;
    assign module_intf_350.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9264.ap_ready;
    assign module_intf_350.ap_done = 1'b0;
    assign module_intf_350.ap_continue = 1'b0;
    assign module_intf_350.finish = finish;
    csv_file_dump mstatus_csv_dumper_350;
    nodf_module_monitor module_monitor_350;
    nodf_module_intf module_intf_351(clock,reset);
    assign module_intf_351.ap_start = 1'b0;
    assign module_intf_351.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9271.ap_ready;
    assign module_intf_351.ap_done = 1'b0;
    assign module_intf_351.ap_continue = 1'b0;
    assign module_intf_351.finish = finish;
    csv_file_dump mstatus_csv_dumper_351;
    nodf_module_monitor module_monitor_351;
    nodf_module_intf module_intf_352(clock,reset);
    assign module_intf_352.ap_start = 1'b0;
    assign module_intf_352.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9278.ap_ready;
    assign module_intf_352.ap_done = 1'b0;
    assign module_intf_352.ap_continue = 1'b0;
    assign module_intf_352.finish = finish;
    csv_file_dump mstatus_csv_dumper_352;
    nodf_module_monitor module_monitor_352;
    nodf_module_intf module_intf_353(clock,reset);
    assign module_intf_353.ap_start = 1'b0;
    assign module_intf_353.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9285.ap_ready;
    assign module_intf_353.ap_done = 1'b0;
    assign module_intf_353.ap_continue = 1'b0;
    assign module_intf_353.finish = finish;
    csv_file_dump mstatus_csv_dumper_353;
    nodf_module_monitor module_monitor_353;
    nodf_module_intf module_intf_354(clock,reset);
    assign module_intf_354.ap_start = 1'b0;
    assign module_intf_354.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9292.ap_ready;
    assign module_intf_354.ap_done = 1'b0;
    assign module_intf_354.ap_continue = 1'b0;
    assign module_intf_354.finish = finish;
    csv_file_dump mstatus_csv_dumper_354;
    nodf_module_monitor module_monitor_354;
    nodf_module_intf module_intf_355(clock,reset);
    assign module_intf_355.ap_start = 1'b0;
    assign module_intf_355.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9299.ap_ready;
    assign module_intf_355.ap_done = 1'b0;
    assign module_intf_355.ap_continue = 1'b0;
    assign module_intf_355.finish = finish;
    csv_file_dump mstatus_csv_dumper_355;
    nodf_module_monitor module_monitor_355;
    nodf_module_intf module_intf_356(clock,reset);
    assign module_intf_356.ap_start = 1'b0;
    assign module_intf_356.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9306.ap_ready;
    assign module_intf_356.ap_done = 1'b0;
    assign module_intf_356.ap_continue = 1'b0;
    assign module_intf_356.finish = finish;
    csv_file_dump mstatus_csv_dumper_356;
    nodf_module_monitor module_monitor_356;
    nodf_module_intf module_intf_357(clock,reset);
    assign module_intf_357.ap_start = 1'b0;
    assign module_intf_357.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9313.ap_ready;
    assign module_intf_357.ap_done = 1'b0;
    assign module_intf_357.ap_continue = 1'b0;
    assign module_intf_357.finish = finish;
    csv_file_dump mstatus_csv_dumper_357;
    nodf_module_monitor module_monitor_357;
    nodf_module_intf module_intf_358(clock,reset);
    assign module_intf_358.ap_start = 1'b0;
    assign module_intf_358.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9320.ap_ready;
    assign module_intf_358.ap_done = 1'b0;
    assign module_intf_358.ap_continue = 1'b0;
    assign module_intf_358.finish = finish;
    csv_file_dump mstatus_csv_dumper_358;
    nodf_module_monitor module_monitor_358;
    nodf_module_intf module_intf_359(clock,reset);
    assign module_intf_359.ap_start = 1'b0;
    assign module_intf_359.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9327.ap_ready;
    assign module_intf_359.ap_done = 1'b0;
    assign module_intf_359.ap_continue = 1'b0;
    assign module_intf_359.finish = finish;
    csv_file_dump mstatus_csv_dumper_359;
    nodf_module_monitor module_monitor_359;
    nodf_module_intf module_intf_360(clock,reset);
    assign module_intf_360.ap_start = 1'b0;
    assign module_intf_360.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9334.ap_ready;
    assign module_intf_360.ap_done = 1'b0;
    assign module_intf_360.ap_continue = 1'b0;
    assign module_intf_360.finish = finish;
    csv_file_dump mstatus_csv_dumper_360;
    nodf_module_monitor module_monitor_360;
    nodf_module_intf module_intf_361(clock,reset);
    assign module_intf_361.ap_start = 1'b0;
    assign module_intf_361.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9341.ap_ready;
    assign module_intf_361.ap_done = 1'b0;
    assign module_intf_361.ap_continue = 1'b0;
    assign module_intf_361.finish = finish;
    csv_file_dump mstatus_csv_dumper_361;
    nodf_module_monitor module_monitor_361;
    nodf_module_intf module_intf_362(clock,reset);
    assign module_intf_362.ap_start = 1'b0;
    assign module_intf_362.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9348.ap_ready;
    assign module_intf_362.ap_done = 1'b0;
    assign module_intf_362.ap_continue = 1'b0;
    assign module_intf_362.finish = finish;
    csv_file_dump mstatus_csv_dumper_362;
    nodf_module_monitor module_monitor_362;
    nodf_module_intf module_intf_363(clock,reset);
    assign module_intf_363.ap_start = 1'b0;
    assign module_intf_363.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9355.ap_ready;
    assign module_intf_363.ap_done = 1'b0;
    assign module_intf_363.ap_continue = 1'b0;
    assign module_intf_363.finish = finish;
    csv_file_dump mstatus_csv_dumper_363;
    nodf_module_monitor module_monitor_363;
    nodf_module_intf module_intf_364(clock,reset);
    assign module_intf_364.ap_start = 1'b0;
    assign module_intf_364.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9362.ap_ready;
    assign module_intf_364.ap_done = 1'b0;
    assign module_intf_364.ap_continue = 1'b0;
    assign module_intf_364.finish = finish;
    csv_file_dump mstatus_csv_dumper_364;
    nodf_module_monitor module_monitor_364;
    nodf_module_intf module_intf_365(clock,reset);
    assign module_intf_365.ap_start = 1'b0;
    assign module_intf_365.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9369.ap_ready;
    assign module_intf_365.ap_done = 1'b0;
    assign module_intf_365.ap_continue = 1'b0;
    assign module_intf_365.finish = finish;
    csv_file_dump mstatus_csv_dumper_365;
    nodf_module_monitor module_monitor_365;
    nodf_module_intf module_intf_366(clock,reset);
    assign module_intf_366.ap_start = 1'b0;
    assign module_intf_366.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9376.ap_ready;
    assign module_intf_366.ap_done = 1'b0;
    assign module_intf_366.ap_continue = 1'b0;
    assign module_intf_366.finish = finish;
    csv_file_dump mstatus_csv_dumper_366;
    nodf_module_monitor module_monitor_366;
    nodf_module_intf module_intf_367(clock,reset);
    assign module_intf_367.ap_start = 1'b0;
    assign module_intf_367.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9383.ap_ready;
    assign module_intf_367.ap_done = 1'b0;
    assign module_intf_367.ap_continue = 1'b0;
    assign module_intf_367.finish = finish;
    csv_file_dump mstatus_csv_dumper_367;
    nodf_module_monitor module_monitor_367;
    nodf_module_intf module_intf_368(clock,reset);
    assign module_intf_368.ap_start = 1'b0;
    assign module_intf_368.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9390.ap_ready;
    assign module_intf_368.ap_done = 1'b0;
    assign module_intf_368.ap_continue = 1'b0;
    assign module_intf_368.finish = finish;
    csv_file_dump mstatus_csv_dumper_368;
    nodf_module_monitor module_monitor_368;
    nodf_module_intf module_intf_369(clock,reset);
    assign module_intf_369.ap_start = 1'b0;
    assign module_intf_369.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9397.ap_ready;
    assign module_intf_369.ap_done = 1'b0;
    assign module_intf_369.ap_continue = 1'b0;
    assign module_intf_369.finish = finish;
    csv_file_dump mstatus_csv_dumper_369;
    nodf_module_monitor module_monitor_369;
    nodf_module_intf module_intf_370(clock,reset);
    assign module_intf_370.ap_start = 1'b0;
    assign module_intf_370.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9404.ap_ready;
    assign module_intf_370.ap_done = 1'b0;
    assign module_intf_370.ap_continue = 1'b0;
    assign module_intf_370.finish = finish;
    csv_file_dump mstatus_csv_dumper_370;
    nodf_module_monitor module_monitor_370;
    nodf_module_intf module_intf_371(clock,reset);
    assign module_intf_371.ap_start = 1'b0;
    assign module_intf_371.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9411.ap_ready;
    assign module_intf_371.ap_done = 1'b0;
    assign module_intf_371.ap_continue = 1'b0;
    assign module_intf_371.finish = finish;
    csv_file_dump mstatus_csv_dumper_371;
    nodf_module_monitor module_monitor_371;
    nodf_module_intf module_intf_372(clock,reset);
    assign module_intf_372.ap_start = 1'b0;
    assign module_intf_372.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9418.ap_ready;
    assign module_intf_372.ap_done = 1'b0;
    assign module_intf_372.ap_continue = 1'b0;
    assign module_intf_372.finish = finish;
    csv_file_dump mstatus_csv_dumper_372;
    nodf_module_monitor module_monitor_372;
    nodf_module_intf module_intf_373(clock,reset);
    assign module_intf_373.ap_start = 1'b0;
    assign module_intf_373.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9425.ap_ready;
    assign module_intf_373.ap_done = 1'b0;
    assign module_intf_373.ap_continue = 1'b0;
    assign module_intf_373.finish = finish;
    csv_file_dump mstatus_csv_dumper_373;
    nodf_module_monitor module_monitor_373;
    nodf_module_intf module_intf_374(clock,reset);
    assign module_intf_374.ap_start = 1'b0;
    assign module_intf_374.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9432.ap_ready;
    assign module_intf_374.ap_done = 1'b0;
    assign module_intf_374.ap_continue = 1'b0;
    assign module_intf_374.finish = finish;
    csv_file_dump mstatus_csv_dumper_374;
    nodf_module_monitor module_monitor_374;
    nodf_module_intf module_intf_375(clock,reset);
    assign module_intf_375.ap_start = 1'b0;
    assign module_intf_375.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9439.ap_ready;
    assign module_intf_375.ap_done = 1'b0;
    assign module_intf_375.ap_continue = 1'b0;
    assign module_intf_375.finish = finish;
    csv_file_dump mstatus_csv_dumper_375;
    nodf_module_monitor module_monitor_375;
    nodf_module_intf module_intf_376(clock,reset);
    assign module_intf_376.ap_start = 1'b0;
    assign module_intf_376.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9446.ap_ready;
    assign module_intf_376.ap_done = 1'b0;
    assign module_intf_376.ap_continue = 1'b0;
    assign module_intf_376.finish = finish;
    csv_file_dump mstatus_csv_dumper_376;
    nodf_module_monitor module_monitor_376;
    nodf_module_intf module_intf_377(clock,reset);
    assign module_intf_377.ap_start = 1'b0;
    assign module_intf_377.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9453.ap_ready;
    assign module_intf_377.ap_done = 1'b0;
    assign module_intf_377.ap_continue = 1'b0;
    assign module_intf_377.finish = finish;
    csv_file_dump mstatus_csv_dumper_377;
    nodf_module_monitor module_monitor_377;
    nodf_module_intf module_intf_378(clock,reset);
    assign module_intf_378.ap_start = 1'b0;
    assign module_intf_378.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9460.ap_ready;
    assign module_intf_378.ap_done = 1'b0;
    assign module_intf_378.ap_continue = 1'b0;
    assign module_intf_378.finish = finish;
    csv_file_dump mstatus_csv_dumper_378;
    nodf_module_monitor module_monitor_378;
    nodf_module_intf module_intf_379(clock,reset);
    assign module_intf_379.ap_start = 1'b0;
    assign module_intf_379.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_add_patch_fu_28570.grp_encodeCoordinates_fu_9467.ap_ready;
    assign module_intf_379.ap_done = 1'b0;
    assign module_intf_379.ap_continue = 1'b0;
    assign module_intf_379.finish = finish;
    csv_file_dump mstatus_csv_dumper_379;
    nodf_module_monitor module_monitor_379;
    nodf_module_intf module_intf_380(clock,reset);
    assign module_intf_380.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.ap_start;
    assign module_intf_380.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.ap_ready;
    assign module_intf_380.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.ap_done;
    assign module_intf_380.ap_continue = 1'b1;
    assign module_intf_380.finish = finish;
    csv_file_dump mstatus_csv_dumper_380;
    nodf_module_monitor module_monitor_380;
    nodf_module_intf module_intf_381(clock,reset);
    assign module_intf_381.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_start;
    assign module_intf_381.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_ready;
    assign module_intf_381.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_done;
    assign module_intf_381.ap_continue = 1'b1;
    assign module_intf_381.finish = finish;
    csv_file_dump mstatus_csv_dumper_381;
    nodf_module_monitor module_monitor_381;
    nodf_module_intf module_intf_382(clock,reset);
    assign module_intf_382.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_start;
    assign module_intf_382.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_ready;
    assign module_intf_382.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_done;
    assign module_intf_382.ap_continue = 1'b1;
    assign module_intf_382.finish = finish;
    csv_file_dump mstatus_csv_dumper_382;
    nodf_module_monitor module_monitor_382;
    nodf_module_intf module_intf_383(clock,reset);
    assign module_intf_383.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_start;
    assign module_intf_383.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_ready;
    assign module_intf_383.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_done;
    assign module_intf_383.ap_continue = 1'b1;
    assign module_intf_383.finish = finish;
    csv_file_dump mstatus_csv_dumper_383;
    nodf_module_monitor module_monitor_383;
    nodf_module_intf module_intf_384(clock,reset);
    assign module_intf_384.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_start;
    assign module_intf_384.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_ready;
    assign module_intf_384.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_done;
    assign module_intf_384.ap_continue = 1'b1;
    assign module_intf_384.finish = finish;
    csv_file_dump mstatus_csv_dumper_384;
    nodf_module_monitor module_monitor_384;
    nodf_module_intf module_intf_385(clock,reset);
    assign module_intf_385.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_start;
    assign module_intf_385.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_ready;
    assign module_intf_385.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_makePatch_alignedToLine_1_fu_48674.grp_wedgePatch_init_fu_29554.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_done;
    assign module_intf_385.ap_continue = 1'b1;
    assign module_intf_385.finish = finish;
    csv_file_dump mstatus_csv_dumper_385;
    nodf_module_monitor module_monitor_385;
    nodf_module_intf module_intf_386(clock,reset);
    assign module_intf_386.ap_start = 1'b0;
    assign module_intf_386.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.tmp_areWedgeSuperPointsEqual_fu_51569.ap_ready;
    assign module_intf_386.ap_done = 1'b0;
    assign module_intf_386.ap_continue = 1'b0;
    assign module_intf_386.finish = finish;
    csv_file_dump mstatus_csv_dumper_386;
    nodf_module_monitor module_monitor_386;
    nodf_module_intf module_intf_387(clock,reset);
    assign module_intf_387.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_straightLineProjectorFromLayerIJtoK_fu_51737.ap_start;
    assign module_intf_387.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_straightLineProjectorFromLayerIJtoK_fu_51737.ap_ready;
    assign module_intf_387.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_straightLineProjectorFromLayerIJtoK_fu_51737.ap_done;
    assign module_intf_387.ap_continue = 1'b1;
    assign module_intf_387.finish = finish;
    csv_file_dump mstatus_csv_dumper_387;
    nodf_module_monitor module_monitor_387;
    nodf_module_intf module_intf_388(clock,reset);
    assign module_intf_388.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_getSolveNextPatchPairWhileCondition_fu_51753.ap_start;
    assign module_intf_388.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_getSolveNextPatchPairWhileCondition_fu_51753.ap_ready;
    assign module_intf_388.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_getSolveNextPatchPairWhileCondition_fu_51753.ap_done;
    assign module_intf_388.ap_continue = 1'b1;
    assign module_intf_388.finish = finish;
    csv_file_dump mstatus_csv_dumper_388;
    nodf_module_monitor module_monitor_388;
    nodf_module_intf module_intf_389(clock,reset);
    assign module_intf_389.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.ap_start;
    assign module_intf_389.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.ap_ready;
    assign module_intf_389.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.ap_done;
    assign module_intf_389.ap_continue = 1'b1;
    assign module_intf_389.finish = finish;
    csv_file_dump mstatus_csv_dumper_389;
    nodf_module_monitor module_monitor_389;
    nodf_module_intf module_intf_390(clock,reset);
    assign module_intf_390.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_start;
    assign module_intf_390.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_ready;
    assign module_intf_390.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.ap_done;
    assign module_intf_390.ap_continue = 1'b1;
    assign module_intf_390.finish = finish;
    csv_file_dump mstatus_csv_dumper_390;
    nodf_module_monitor module_monitor_390;
    nodf_module_intf module_intf_391(clock,reset);
    assign module_intf_391.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_start;
    assign module_intf_391.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_ready;
    assign module_intf_391.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_322.ap_done;
    assign module_intf_391.ap_continue = 1'b1;
    assign module_intf_391.finish = finish;
    csv_file_dump mstatus_csv_dumper_391;
    nodf_module_monitor module_monitor_391;
    nodf_module_intf module_intf_392(clock,reset);
    assign module_intf_392.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_start;
    assign module_intf_392.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_ready;
    assign module_intf_392.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_335.ap_done;
    assign module_intf_392.ap_continue = 1'b1;
    assign module_intf_392.finish = finish;
    csv_file_dump mstatus_csv_dumper_392;
    nodf_module_monitor module_monitor_392;
    nodf_module_intf module_intf_393(clock,reset);
    assign module_intf_393.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_start;
    assign module_intf_393.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_ready;
    assign module_intf_393.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_348.ap_done;
    assign module_intf_393.ap_continue = 1'b1;
    assign module_intf_393.finish = finish;
    csv_file_dump mstatus_csv_dumper_393;
    nodf_module_monitor module_monitor_393;
    nodf_module_intf module_intf_394(clock,reset);
    assign module_intf_394.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_start;
    assign module_intf_394.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_ready;
    assign module_intf_394.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_wedgePatch_init_fu_86940.grp_getParallelogramsAndAcceptanceCorners_fu_2673.grp_straightLineProjectorFromLayerIJtoK_fu_362.ap_done;
    assign module_intf_394.ap_continue = 1'b1;
    assign module_intf_394.finish = finish;
    csv_file_dump mstatus_csv_dumper_394;
    nodf_module_monitor module_monitor_394;
    nodf_module_intf module_intf_395(clock,reset);
    assign module_intf_395.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_straightLineProjectorFromLayerIJtoK_fu_87108.ap_start;
    assign module_intf_395.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_straightLineProjectorFromLayerIJtoK_fu_87108.ap_ready;
    assign module_intf_395.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_solveNextPatchPair_fu_29444.grp_straightLineProjectorFromLayerIJtoK_fu_87108.ap_done;
    assign module_intf_395.ap_continue = 1'b1;
    assign module_intf_395.finish = finish;
    csv_file_dump mstatus_csv_dumper_395;
    nodf_module_monitor module_monitor_395;
    nodf_module_intf module_intf_396(clock,reset);
    assign module_intf_396.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_straightLineProjectorFromLayerIJtoK_fu_32657.ap_start;
    assign module_intf_396.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_straightLineProjectorFromLayerIJtoK_fu_32657.ap_ready;
    assign module_intf_396.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.grp_straightLineProjectorFromLayerIJtoK_fu_32657.ap_done;
    assign module_intf_396.ap_continue = 1'b1;
    assign module_intf_396.finish = finish;
    csv_file_dump mstatus_csv_dumper_396;
    nodf_module_monitor module_monitor_396;
    nodf_module_intf module_intf_397(clock,reset);
    assign module_intf_397.ap_start = 1'b0;
    assign module_intf_397.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_20111.tmp_getSolveNextColumnWhileConditional_fu_32673.ap_ready;
    assign module_intf_397.ap_done = 1'b0;
    assign module_intf_397.ap_continue = 1'b0;
    assign module_intf_397.finish = finish;
    csv_file_dump mstatus_csv_dumper_397;
    nodf_module_monitor module_monitor_397;
    nodf_module_intf module_intf_398(clock,reset);
    assign module_intf_398.ap_start = AESL_inst_MPSQ.grp_initializeArrays_fu_23317.ap_start;
    assign module_intf_398.ap_ready = AESL_inst_MPSQ.grp_initializeArrays_fu_23317.ap_ready;
    assign module_intf_398.ap_done = AESL_inst_MPSQ.grp_initializeArrays_fu_23317.ap_done;
    assign module_intf_398.ap_continue = 1'b1;
    assign module_intf_398.finish = finish;
    csv_file_dump mstatus_csv_dumper_398;
    nodf_module_monitor module_monitor_398;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);
    mstatus_csv_dumper_58 = new("./module_status58.csv");
    module_monitor_58 = new(module_intf_58,mstatus_csv_dumper_58);
    mstatus_csv_dumper_59 = new("./module_status59.csv");
    module_monitor_59 = new(module_intf_59,mstatus_csv_dumper_59);
    mstatus_csv_dumper_60 = new("./module_status60.csv");
    module_monitor_60 = new(module_intf_60,mstatus_csv_dumper_60);
    mstatus_csv_dumper_61 = new("./module_status61.csv");
    module_monitor_61 = new(module_intf_61,mstatus_csv_dumper_61);
    mstatus_csv_dumper_62 = new("./module_status62.csv");
    module_monitor_62 = new(module_intf_62,mstatus_csv_dumper_62);
    mstatus_csv_dumper_63 = new("./module_status63.csv");
    module_monitor_63 = new(module_intf_63,mstatus_csv_dumper_63);
    mstatus_csv_dumper_64 = new("./module_status64.csv");
    module_monitor_64 = new(module_intf_64,mstatus_csv_dumper_64);
    mstatus_csv_dumper_65 = new("./module_status65.csv");
    module_monitor_65 = new(module_intf_65,mstatus_csv_dumper_65);
    mstatus_csv_dumper_66 = new("./module_status66.csv");
    module_monitor_66 = new(module_intf_66,mstatus_csv_dumper_66);
    mstatus_csv_dumper_67 = new("./module_status67.csv");
    module_monitor_67 = new(module_intf_67,mstatus_csv_dumper_67);
    mstatus_csv_dumper_68 = new("./module_status68.csv");
    module_monitor_68 = new(module_intf_68,mstatus_csv_dumper_68);
    mstatus_csv_dumper_69 = new("./module_status69.csv");
    module_monitor_69 = new(module_intf_69,mstatus_csv_dumper_69);
    mstatus_csv_dumper_70 = new("./module_status70.csv");
    module_monitor_70 = new(module_intf_70,mstatus_csv_dumper_70);
    mstatus_csv_dumper_71 = new("./module_status71.csv");
    module_monitor_71 = new(module_intf_71,mstatus_csv_dumper_71);
    mstatus_csv_dumper_72 = new("./module_status72.csv");
    module_monitor_72 = new(module_intf_72,mstatus_csv_dumper_72);
    mstatus_csv_dumper_73 = new("./module_status73.csv");
    module_monitor_73 = new(module_intf_73,mstatus_csv_dumper_73);
    mstatus_csv_dumper_74 = new("./module_status74.csv");
    module_monitor_74 = new(module_intf_74,mstatus_csv_dumper_74);
    mstatus_csv_dumper_75 = new("./module_status75.csv");
    module_monitor_75 = new(module_intf_75,mstatus_csv_dumper_75);
    mstatus_csv_dumper_76 = new("./module_status76.csv");
    module_monitor_76 = new(module_intf_76,mstatus_csv_dumper_76);
    mstatus_csv_dumper_77 = new("./module_status77.csv");
    module_monitor_77 = new(module_intf_77,mstatus_csv_dumper_77);
    mstatus_csv_dumper_78 = new("./module_status78.csv");
    module_monitor_78 = new(module_intf_78,mstatus_csv_dumper_78);
    mstatus_csv_dumper_79 = new("./module_status79.csv");
    module_monitor_79 = new(module_intf_79,mstatus_csv_dumper_79);
    mstatus_csv_dumper_80 = new("./module_status80.csv");
    module_monitor_80 = new(module_intf_80,mstatus_csv_dumper_80);
    mstatus_csv_dumper_81 = new("./module_status81.csv");
    module_monitor_81 = new(module_intf_81,mstatus_csv_dumper_81);
    mstatus_csv_dumper_82 = new("./module_status82.csv");
    module_monitor_82 = new(module_intf_82,mstatus_csv_dumper_82);
    mstatus_csv_dumper_83 = new("./module_status83.csv");
    module_monitor_83 = new(module_intf_83,mstatus_csv_dumper_83);
    mstatus_csv_dumper_84 = new("./module_status84.csv");
    module_monitor_84 = new(module_intf_84,mstatus_csv_dumper_84);
    mstatus_csv_dumper_85 = new("./module_status85.csv");
    module_monitor_85 = new(module_intf_85,mstatus_csv_dumper_85);
    mstatus_csv_dumper_86 = new("./module_status86.csv");
    module_monitor_86 = new(module_intf_86,mstatus_csv_dumper_86);
    mstatus_csv_dumper_87 = new("./module_status87.csv");
    module_monitor_87 = new(module_intf_87,mstatus_csv_dumper_87);
    mstatus_csv_dumper_88 = new("./module_status88.csv");
    module_monitor_88 = new(module_intf_88,mstatus_csv_dumper_88);
    mstatus_csv_dumper_89 = new("./module_status89.csv");
    module_monitor_89 = new(module_intf_89,mstatus_csv_dumper_89);
    mstatus_csv_dumper_90 = new("./module_status90.csv");
    module_monitor_90 = new(module_intf_90,mstatus_csv_dumper_90);
    mstatus_csv_dumper_91 = new("./module_status91.csv");
    module_monitor_91 = new(module_intf_91,mstatus_csv_dumper_91);
    mstatus_csv_dumper_92 = new("./module_status92.csv");
    module_monitor_92 = new(module_intf_92,mstatus_csv_dumper_92);
    mstatus_csv_dumper_93 = new("./module_status93.csv");
    module_monitor_93 = new(module_intf_93,mstatus_csv_dumper_93);
    mstatus_csv_dumper_94 = new("./module_status94.csv");
    module_monitor_94 = new(module_intf_94,mstatus_csv_dumper_94);
    mstatus_csv_dumper_95 = new("./module_status95.csv");
    module_monitor_95 = new(module_intf_95,mstatus_csv_dumper_95);
    mstatus_csv_dumper_96 = new("./module_status96.csv");
    module_monitor_96 = new(module_intf_96,mstatus_csv_dumper_96);
    mstatus_csv_dumper_97 = new("./module_status97.csv");
    module_monitor_97 = new(module_intf_97,mstatus_csv_dumper_97);
    mstatus_csv_dumper_98 = new("./module_status98.csv");
    module_monitor_98 = new(module_intf_98,mstatus_csv_dumper_98);
    mstatus_csv_dumper_99 = new("./module_status99.csv");
    module_monitor_99 = new(module_intf_99,mstatus_csv_dumper_99);
    mstatus_csv_dumper_100 = new("./module_status100.csv");
    module_monitor_100 = new(module_intf_100,mstatus_csv_dumper_100);
    mstatus_csv_dumper_101 = new("./module_status101.csv");
    module_monitor_101 = new(module_intf_101,mstatus_csv_dumper_101);
    mstatus_csv_dumper_102 = new("./module_status102.csv");
    module_monitor_102 = new(module_intf_102,mstatus_csv_dumper_102);
    mstatus_csv_dumper_103 = new("./module_status103.csv");
    module_monitor_103 = new(module_intf_103,mstatus_csv_dumper_103);
    mstatus_csv_dumper_104 = new("./module_status104.csv");
    module_monitor_104 = new(module_intf_104,mstatus_csv_dumper_104);
    mstatus_csv_dumper_105 = new("./module_status105.csv");
    module_monitor_105 = new(module_intf_105,mstatus_csv_dumper_105);
    mstatus_csv_dumper_106 = new("./module_status106.csv");
    module_monitor_106 = new(module_intf_106,mstatus_csv_dumper_106);
    mstatus_csv_dumper_107 = new("./module_status107.csv");
    module_monitor_107 = new(module_intf_107,mstatus_csv_dumper_107);
    mstatus_csv_dumper_108 = new("./module_status108.csv");
    module_monitor_108 = new(module_intf_108,mstatus_csv_dumper_108);
    mstatus_csv_dumper_109 = new("./module_status109.csv");
    module_monitor_109 = new(module_intf_109,mstatus_csv_dumper_109);
    mstatus_csv_dumper_110 = new("./module_status110.csv");
    module_monitor_110 = new(module_intf_110,mstatus_csv_dumper_110);
    mstatus_csv_dumper_111 = new("./module_status111.csv");
    module_monitor_111 = new(module_intf_111,mstatus_csv_dumper_111);
    mstatus_csv_dumper_112 = new("./module_status112.csv");
    module_monitor_112 = new(module_intf_112,mstatus_csv_dumper_112);
    mstatus_csv_dumper_113 = new("./module_status113.csv");
    module_monitor_113 = new(module_intf_113,mstatus_csv_dumper_113);
    mstatus_csv_dumper_114 = new("./module_status114.csv");
    module_monitor_114 = new(module_intf_114,mstatus_csv_dumper_114);
    mstatus_csv_dumper_115 = new("./module_status115.csv");
    module_monitor_115 = new(module_intf_115,mstatus_csv_dumper_115);
    mstatus_csv_dumper_116 = new("./module_status116.csv");
    module_monitor_116 = new(module_intf_116,mstatus_csv_dumper_116);
    mstatus_csv_dumper_117 = new("./module_status117.csv");
    module_monitor_117 = new(module_intf_117,mstatus_csv_dumper_117);
    mstatus_csv_dumper_118 = new("./module_status118.csv");
    module_monitor_118 = new(module_intf_118,mstatus_csv_dumper_118);
    mstatus_csv_dumper_119 = new("./module_status119.csv");
    module_monitor_119 = new(module_intf_119,mstatus_csv_dumper_119);
    mstatus_csv_dumper_120 = new("./module_status120.csv");
    module_monitor_120 = new(module_intf_120,mstatus_csv_dumper_120);
    mstatus_csv_dumper_121 = new("./module_status121.csv");
    module_monitor_121 = new(module_intf_121,mstatus_csv_dumper_121);
    mstatus_csv_dumper_122 = new("./module_status122.csv");
    module_monitor_122 = new(module_intf_122,mstatus_csv_dumper_122);
    mstatus_csv_dumper_123 = new("./module_status123.csv");
    module_monitor_123 = new(module_intf_123,mstatus_csv_dumper_123);
    mstatus_csv_dumper_124 = new("./module_status124.csv");
    module_monitor_124 = new(module_intf_124,mstatus_csv_dumper_124);
    mstatus_csv_dumper_125 = new("./module_status125.csv");
    module_monitor_125 = new(module_intf_125,mstatus_csv_dumper_125);
    mstatus_csv_dumper_126 = new("./module_status126.csv");
    module_monitor_126 = new(module_intf_126,mstatus_csv_dumper_126);
    mstatus_csv_dumper_127 = new("./module_status127.csv");
    module_monitor_127 = new(module_intf_127,mstatus_csv_dumper_127);
    mstatus_csv_dumper_128 = new("./module_status128.csv");
    module_monitor_128 = new(module_intf_128,mstatus_csv_dumper_128);
    mstatus_csv_dumper_129 = new("./module_status129.csv");
    module_monitor_129 = new(module_intf_129,mstatus_csv_dumper_129);
    mstatus_csv_dumper_130 = new("./module_status130.csv");
    module_monitor_130 = new(module_intf_130,mstatus_csv_dumper_130);
    mstatus_csv_dumper_131 = new("./module_status131.csv");
    module_monitor_131 = new(module_intf_131,mstatus_csv_dumper_131);
    mstatus_csv_dumper_132 = new("./module_status132.csv");
    module_monitor_132 = new(module_intf_132,mstatus_csv_dumper_132);
    mstatus_csv_dumper_133 = new("./module_status133.csv");
    module_monitor_133 = new(module_intf_133,mstatus_csv_dumper_133);
    mstatus_csv_dumper_134 = new("./module_status134.csv");
    module_monitor_134 = new(module_intf_134,mstatus_csv_dumper_134);
    mstatus_csv_dumper_135 = new("./module_status135.csv");
    module_monitor_135 = new(module_intf_135,mstatus_csv_dumper_135);
    mstatus_csv_dumper_136 = new("./module_status136.csv");
    module_monitor_136 = new(module_intf_136,mstatus_csv_dumper_136);
    mstatus_csv_dumper_137 = new("./module_status137.csv");
    module_monitor_137 = new(module_intf_137,mstatus_csv_dumper_137);
    mstatus_csv_dumper_138 = new("./module_status138.csv");
    module_monitor_138 = new(module_intf_138,mstatus_csv_dumper_138);
    mstatus_csv_dumper_139 = new("./module_status139.csv");
    module_monitor_139 = new(module_intf_139,mstatus_csv_dumper_139);
    mstatus_csv_dumper_140 = new("./module_status140.csv");
    module_monitor_140 = new(module_intf_140,mstatus_csv_dumper_140);
    mstatus_csv_dumper_141 = new("./module_status141.csv");
    module_monitor_141 = new(module_intf_141,mstatus_csv_dumper_141);
    mstatus_csv_dumper_142 = new("./module_status142.csv");
    module_monitor_142 = new(module_intf_142,mstatus_csv_dumper_142);
    mstatus_csv_dumper_143 = new("./module_status143.csv");
    module_monitor_143 = new(module_intf_143,mstatus_csv_dumper_143);
    mstatus_csv_dumper_144 = new("./module_status144.csv");
    module_monitor_144 = new(module_intf_144,mstatus_csv_dumper_144);
    mstatus_csv_dumper_145 = new("./module_status145.csv");
    module_monitor_145 = new(module_intf_145,mstatus_csv_dumper_145);
    mstatus_csv_dumper_146 = new("./module_status146.csv");
    module_monitor_146 = new(module_intf_146,mstatus_csv_dumper_146);
    mstatus_csv_dumper_147 = new("./module_status147.csv");
    module_monitor_147 = new(module_intf_147,mstatus_csv_dumper_147);
    mstatus_csv_dumper_148 = new("./module_status148.csv");
    module_monitor_148 = new(module_intf_148,mstatus_csv_dumper_148);
    mstatus_csv_dumper_149 = new("./module_status149.csv");
    module_monitor_149 = new(module_intf_149,mstatus_csv_dumper_149);
    mstatus_csv_dumper_150 = new("./module_status150.csv");
    module_monitor_150 = new(module_intf_150,mstatus_csv_dumper_150);
    mstatus_csv_dumper_151 = new("./module_status151.csv");
    module_monitor_151 = new(module_intf_151,mstatus_csv_dumper_151);
    mstatus_csv_dumper_152 = new("./module_status152.csv");
    module_monitor_152 = new(module_intf_152,mstatus_csv_dumper_152);
    mstatus_csv_dumper_153 = new("./module_status153.csv");
    module_monitor_153 = new(module_intf_153,mstatus_csv_dumper_153);
    mstatus_csv_dumper_154 = new("./module_status154.csv");
    module_monitor_154 = new(module_intf_154,mstatus_csv_dumper_154);
    mstatus_csv_dumper_155 = new("./module_status155.csv");
    module_monitor_155 = new(module_intf_155,mstatus_csv_dumper_155);
    mstatus_csv_dumper_156 = new("./module_status156.csv");
    module_monitor_156 = new(module_intf_156,mstatus_csv_dumper_156);
    mstatus_csv_dumper_157 = new("./module_status157.csv");
    module_monitor_157 = new(module_intf_157,mstatus_csv_dumper_157);
    mstatus_csv_dumper_158 = new("./module_status158.csv");
    module_monitor_158 = new(module_intf_158,mstatus_csv_dumper_158);
    mstatus_csv_dumper_159 = new("./module_status159.csv");
    module_monitor_159 = new(module_intf_159,mstatus_csv_dumper_159);
    mstatus_csv_dumper_160 = new("./module_status160.csv");
    module_monitor_160 = new(module_intf_160,mstatus_csv_dumper_160);
    mstatus_csv_dumper_161 = new("./module_status161.csv");
    module_monitor_161 = new(module_intf_161,mstatus_csv_dumper_161);
    mstatus_csv_dumper_162 = new("./module_status162.csv");
    module_monitor_162 = new(module_intf_162,mstatus_csv_dumper_162);
    mstatus_csv_dumper_163 = new("./module_status163.csv");
    module_monitor_163 = new(module_intf_163,mstatus_csv_dumper_163);
    mstatus_csv_dumper_164 = new("./module_status164.csv");
    module_monitor_164 = new(module_intf_164,mstatus_csv_dumper_164);
    mstatus_csv_dumper_165 = new("./module_status165.csv");
    module_monitor_165 = new(module_intf_165,mstatus_csv_dumper_165);
    mstatus_csv_dumper_166 = new("./module_status166.csv");
    module_monitor_166 = new(module_intf_166,mstatus_csv_dumper_166);
    mstatus_csv_dumper_167 = new("./module_status167.csv");
    module_monitor_167 = new(module_intf_167,mstatus_csv_dumper_167);
    mstatus_csv_dumper_168 = new("./module_status168.csv");
    module_monitor_168 = new(module_intf_168,mstatus_csv_dumper_168);
    mstatus_csv_dumper_169 = new("./module_status169.csv");
    module_monitor_169 = new(module_intf_169,mstatus_csv_dumper_169);
    mstatus_csv_dumper_170 = new("./module_status170.csv");
    module_monitor_170 = new(module_intf_170,mstatus_csv_dumper_170);
    mstatus_csv_dumper_171 = new("./module_status171.csv");
    module_monitor_171 = new(module_intf_171,mstatus_csv_dumper_171);
    mstatus_csv_dumper_172 = new("./module_status172.csv");
    module_monitor_172 = new(module_intf_172,mstatus_csv_dumper_172);
    mstatus_csv_dumper_173 = new("./module_status173.csv");
    module_monitor_173 = new(module_intf_173,mstatus_csv_dumper_173);
    mstatus_csv_dumper_174 = new("./module_status174.csv");
    module_monitor_174 = new(module_intf_174,mstatus_csv_dumper_174);
    mstatus_csv_dumper_175 = new("./module_status175.csv");
    module_monitor_175 = new(module_intf_175,mstatus_csv_dumper_175);
    mstatus_csv_dumper_176 = new("./module_status176.csv");
    module_monitor_176 = new(module_intf_176,mstatus_csv_dumper_176);
    mstatus_csv_dumper_177 = new("./module_status177.csv");
    module_monitor_177 = new(module_intf_177,mstatus_csv_dumper_177);
    mstatus_csv_dumper_178 = new("./module_status178.csv");
    module_monitor_178 = new(module_intf_178,mstatus_csv_dumper_178);
    mstatus_csv_dumper_179 = new("./module_status179.csv");
    module_monitor_179 = new(module_intf_179,mstatus_csv_dumper_179);
    mstatus_csv_dumper_180 = new("./module_status180.csv");
    module_monitor_180 = new(module_intf_180,mstatus_csv_dumper_180);
    mstatus_csv_dumper_181 = new("./module_status181.csv");
    module_monitor_181 = new(module_intf_181,mstatus_csv_dumper_181);
    mstatus_csv_dumper_182 = new("./module_status182.csv");
    module_monitor_182 = new(module_intf_182,mstatus_csv_dumper_182);
    mstatus_csv_dumper_183 = new("./module_status183.csv");
    module_monitor_183 = new(module_intf_183,mstatus_csv_dumper_183);
    mstatus_csv_dumper_184 = new("./module_status184.csv");
    module_monitor_184 = new(module_intf_184,mstatus_csv_dumper_184);
    mstatus_csv_dumper_185 = new("./module_status185.csv");
    module_monitor_185 = new(module_intf_185,mstatus_csv_dumper_185);
    mstatus_csv_dumper_186 = new("./module_status186.csv");
    module_monitor_186 = new(module_intf_186,mstatus_csv_dumper_186);
    mstatus_csv_dumper_187 = new("./module_status187.csv");
    module_monitor_187 = new(module_intf_187,mstatus_csv_dumper_187);
    mstatus_csv_dumper_188 = new("./module_status188.csv");
    module_monitor_188 = new(module_intf_188,mstatus_csv_dumper_188);
    mstatus_csv_dumper_189 = new("./module_status189.csv");
    module_monitor_189 = new(module_intf_189,mstatus_csv_dumper_189);
    mstatus_csv_dumper_190 = new("./module_status190.csv");
    module_monitor_190 = new(module_intf_190,mstatus_csv_dumper_190);
    mstatus_csv_dumper_191 = new("./module_status191.csv");
    module_monitor_191 = new(module_intf_191,mstatus_csv_dumper_191);
    mstatus_csv_dumper_192 = new("./module_status192.csv");
    module_monitor_192 = new(module_intf_192,mstatus_csv_dumper_192);
    mstatus_csv_dumper_193 = new("./module_status193.csv");
    module_monitor_193 = new(module_intf_193,mstatus_csv_dumper_193);
    mstatus_csv_dumper_194 = new("./module_status194.csv");
    module_monitor_194 = new(module_intf_194,mstatus_csv_dumper_194);
    mstatus_csv_dumper_195 = new("./module_status195.csv");
    module_monitor_195 = new(module_intf_195,mstatus_csv_dumper_195);
    mstatus_csv_dumper_196 = new("./module_status196.csv");
    module_monitor_196 = new(module_intf_196,mstatus_csv_dumper_196);
    mstatus_csv_dumper_197 = new("./module_status197.csv");
    module_monitor_197 = new(module_intf_197,mstatus_csv_dumper_197);
    mstatus_csv_dumper_198 = new("./module_status198.csv");
    module_monitor_198 = new(module_intf_198,mstatus_csv_dumper_198);
    mstatus_csv_dumper_199 = new("./module_status199.csv");
    module_monitor_199 = new(module_intf_199,mstatus_csv_dumper_199);
    mstatus_csv_dumper_200 = new("./module_status200.csv");
    module_monitor_200 = new(module_intf_200,mstatus_csv_dumper_200);
    mstatus_csv_dumper_201 = new("./module_status201.csv");
    module_monitor_201 = new(module_intf_201,mstatus_csv_dumper_201);
    mstatus_csv_dumper_202 = new("./module_status202.csv");
    module_monitor_202 = new(module_intf_202,mstatus_csv_dumper_202);
    mstatus_csv_dumper_203 = new("./module_status203.csv");
    module_monitor_203 = new(module_intf_203,mstatus_csv_dumper_203);
    mstatus_csv_dumper_204 = new("./module_status204.csv");
    module_monitor_204 = new(module_intf_204,mstatus_csv_dumper_204);
    mstatus_csv_dumper_205 = new("./module_status205.csv");
    module_monitor_205 = new(module_intf_205,mstatus_csv_dumper_205);
    mstatus_csv_dumper_206 = new("./module_status206.csv");
    module_monitor_206 = new(module_intf_206,mstatus_csv_dumper_206);
    mstatus_csv_dumper_207 = new("./module_status207.csv");
    module_monitor_207 = new(module_intf_207,mstatus_csv_dumper_207);
    mstatus_csv_dumper_208 = new("./module_status208.csv");
    module_monitor_208 = new(module_intf_208,mstatus_csv_dumper_208);
    mstatus_csv_dumper_209 = new("./module_status209.csv");
    module_monitor_209 = new(module_intf_209,mstatus_csv_dumper_209);
    mstatus_csv_dumper_210 = new("./module_status210.csv");
    module_monitor_210 = new(module_intf_210,mstatus_csv_dumper_210);
    mstatus_csv_dumper_211 = new("./module_status211.csv");
    module_monitor_211 = new(module_intf_211,mstatus_csv_dumper_211);
    mstatus_csv_dumper_212 = new("./module_status212.csv");
    module_monitor_212 = new(module_intf_212,mstatus_csv_dumper_212);
    mstatus_csv_dumper_213 = new("./module_status213.csv");
    module_monitor_213 = new(module_intf_213,mstatus_csv_dumper_213);
    mstatus_csv_dumper_214 = new("./module_status214.csv");
    module_monitor_214 = new(module_intf_214,mstatus_csv_dumper_214);
    mstatus_csv_dumper_215 = new("./module_status215.csv");
    module_monitor_215 = new(module_intf_215,mstatus_csv_dumper_215);
    mstatus_csv_dumper_216 = new("./module_status216.csv");
    module_monitor_216 = new(module_intf_216,mstatus_csv_dumper_216);
    mstatus_csv_dumper_217 = new("./module_status217.csv");
    module_monitor_217 = new(module_intf_217,mstatus_csv_dumper_217);
    mstatus_csv_dumper_218 = new("./module_status218.csv");
    module_monitor_218 = new(module_intf_218,mstatus_csv_dumper_218);
    mstatus_csv_dumper_219 = new("./module_status219.csv");
    module_monitor_219 = new(module_intf_219,mstatus_csv_dumper_219);
    mstatus_csv_dumper_220 = new("./module_status220.csv");
    module_monitor_220 = new(module_intf_220,mstatus_csv_dumper_220);
    mstatus_csv_dumper_221 = new("./module_status221.csv");
    module_monitor_221 = new(module_intf_221,mstatus_csv_dumper_221);
    mstatus_csv_dumper_222 = new("./module_status222.csv");
    module_monitor_222 = new(module_intf_222,mstatus_csv_dumper_222);
    mstatus_csv_dumper_223 = new("./module_status223.csv");
    module_monitor_223 = new(module_intf_223,mstatus_csv_dumper_223);
    mstatus_csv_dumper_224 = new("./module_status224.csv");
    module_monitor_224 = new(module_intf_224,mstatus_csv_dumper_224);
    mstatus_csv_dumper_225 = new("./module_status225.csv");
    module_monitor_225 = new(module_intf_225,mstatus_csv_dumper_225);
    mstatus_csv_dumper_226 = new("./module_status226.csv");
    module_monitor_226 = new(module_intf_226,mstatus_csv_dumper_226);
    mstatus_csv_dumper_227 = new("./module_status227.csv");
    module_monitor_227 = new(module_intf_227,mstatus_csv_dumper_227);
    mstatus_csv_dumper_228 = new("./module_status228.csv");
    module_monitor_228 = new(module_intf_228,mstatus_csv_dumper_228);
    mstatus_csv_dumper_229 = new("./module_status229.csv");
    module_monitor_229 = new(module_intf_229,mstatus_csv_dumper_229);
    mstatus_csv_dumper_230 = new("./module_status230.csv");
    module_monitor_230 = new(module_intf_230,mstatus_csv_dumper_230);
    mstatus_csv_dumper_231 = new("./module_status231.csv");
    module_monitor_231 = new(module_intf_231,mstatus_csv_dumper_231);
    mstatus_csv_dumper_232 = new("./module_status232.csv");
    module_monitor_232 = new(module_intf_232,mstatus_csv_dumper_232);
    mstatus_csv_dumper_233 = new("./module_status233.csv");
    module_monitor_233 = new(module_intf_233,mstatus_csv_dumper_233);
    mstatus_csv_dumper_234 = new("./module_status234.csv");
    module_monitor_234 = new(module_intf_234,mstatus_csv_dumper_234);
    mstatus_csv_dumper_235 = new("./module_status235.csv");
    module_monitor_235 = new(module_intf_235,mstatus_csv_dumper_235);
    mstatus_csv_dumper_236 = new("./module_status236.csv");
    module_monitor_236 = new(module_intf_236,mstatus_csv_dumper_236);
    mstatus_csv_dumper_237 = new("./module_status237.csv");
    module_monitor_237 = new(module_intf_237,mstatus_csv_dumper_237);
    mstatus_csv_dumper_238 = new("./module_status238.csv");
    module_monitor_238 = new(module_intf_238,mstatus_csv_dumper_238);
    mstatus_csv_dumper_239 = new("./module_status239.csv");
    module_monitor_239 = new(module_intf_239,mstatus_csv_dumper_239);
    mstatus_csv_dumper_240 = new("./module_status240.csv");
    module_monitor_240 = new(module_intf_240,mstatus_csv_dumper_240);
    mstatus_csv_dumper_241 = new("./module_status241.csv");
    module_monitor_241 = new(module_intf_241,mstatus_csv_dumper_241);
    mstatus_csv_dumper_242 = new("./module_status242.csv");
    module_monitor_242 = new(module_intf_242,mstatus_csv_dumper_242);
    mstatus_csv_dumper_243 = new("./module_status243.csv");
    module_monitor_243 = new(module_intf_243,mstatus_csv_dumper_243);
    mstatus_csv_dumper_244 = new("./module_status244.csv");
    module_monitor_244 = new(module_intf_244,mstatus_csv_dumper_244);
    mstatus_csv_dumper_245 = new("./module_status245.csv");
    module_monitor_245 = new(module_intf_245,mstatus_csv_dumper_245);
    mstatus_csv_dumper_246 = new("./module_status246.csv");
    module_monitor_246 = new(module_intf_246,mstatus_csv_dumper_246);
    mstatus_csv_dumper_247 = new("./module_status247.csv");
    module_monitor_247 = new(module_intf_247,mstatus_csv_dumper_247);
    mstatus_csv_dumper_248 = new("./module_status248.csv");
    module_monitor_248 = new(module_intf_248,mstatus_csv_dumper_248);
    mstatus_csv_dumper_249 = new("./module_status249.csv");
    module_monitor_249 = new(module_intf_249,mstatus_csv_dumper_249);
    mstatus_csv_dumper_250 = new("./module_status250.csv");
    module_monitor_250 = new(module_intf_250,mstatus_csv_dumper_250);
    mstatus_csv_dumper_251 = new("./module_status251.csv");
    module_monitor_251 = new(module_intf_251,mstatus_csv_dumper_251);
    mstatus_csv_dumper_252 = new("./module_status252.csv");
    module_monitor_252 = new(module_intf_252,mstatus_csv_dumper_252);
    mstatus_csv_dumper_253 = new("./module_status253.csv");
    module_monitor_253 = new(module_intf_253,mstatus_csv_dumper_253);
    mstatus_csv_dumper_254 = new("./module_status254.csv");
    module_monitor_254 = new(module_intf_254,mstatus_csv_dumper_254);
    mstatus_csv_dumper_255 = new("./module_status255.csv");
    module_monitor_255 = new(module_intf_255,mstatus_csv_dumper_255);
    mstatus_csv_dumper_256 = new("./module_status256.csv");
    module_monitor_256 = new(module_intf_256,mstatus_csv_dumper_256);
    mstatus_csv_dumper_257 = new("./module_status257.csv");
    module_monitor_257 = new(module_intf_257,mstatus_csv_dumper_257);
    mstatus_csv_dumper_258 = new("./module_status258.csv");
    module_monitor_258 = new(module_intf_258,mstatus_csv_dumper_258);
    mstatus_csv_dumper_259 = new("./module_status259.csv");
    module_monitor_259 = new(module_intf_259,mstatus_csv_dumper_259);
    mstatus_csv_dumper_260 = new("./module_status260.csv");
    module_monitor_260 = new(module_intf_260,mstatus_csv_dumper_260);
    mstatus_csv_dumper_261 = new("./module_status261.csv");
    module_monitor_261 = new(module_intf_261,mstatus_csv_dumper_261);
    mstatus_csv_dumper_262 = new("./module_status262.csv");
    module_monitor_262 = new(module_intf_262,mstatus_csv_dumper_262);
    mstatus_csv_dumper_263 = new("./module_status263.csv");
    module_monitor_263 = new(module_intf_263,mstatus_csv_dumper_263);
    mstatus_csv_dumper_264 = new("./module_status264.csv");
    module_monitor_264 = new(module_intf_264,mstatus_csv_dumper_264);
    mstatus_csv_dumper_265 = new("./module_status265.csv");
    module_monitor_265 = new(module_intf_265,mstatus_csv_dumper_265);
    mstatus_csv_dumper_266 = new("./module_status266.csv");
    module_monitor_266 = new(module_intf_266,mstatus_csv_dumper_266);
    mstatus_csv_dumper_267 = new("./module_status267.csv");
    module_monitor_267 = new(module_intf_267,mstatus_csv_dumper_267);
    mstatus_csv_dumper_268 = new("./module_status268.csv");
    module_monitor_268 = new(module_intf_268,mstatus_csv_dumper_268);
    mstatus_csv_dumper_269 = new("./module_status269.csv");
    module_monitor_269 = new(module_intf_269,mstatus_csv_dumper_269);
    mstatus_csv_dumper_270 = new("./module_status270.csv");
    module_monitor_270 = new(module_intf_270,mstatus_csv_dumper_270);
    mstatus_csv_dumper_271 = new("./module_status271.csv");
    module_monitor_271 = new(module_intf_271,mstatus_csv_dumper_271);
    mstatus_csv_dumper_272 = new("./module_status272.csv");
    module_monitor_272 = new(module_intf_272,mstatus_csv_dumper_272);
    mstatus_csv_dumper_273 = new("./module_status273.csv");
    module_monitor_273 = new(module_intf_273,mstatus_csv_dumper_273);
    mstatus_csv_dumper_274 = new("./module_status274.csv");
    module_monitor_274 = new(module_intf_274,mstatus_csv_dumper_274);
    mstatus_csv_dumper_275 = new("./module_status275.csv");
    module_monitor_275 = new(module_intf_275,mstatus_csv_dumper_275);
    mstatus_csv_dumper_276 = new("./module_status276.csv");
    module_monitor_276 = new(module_intf_276,mstatus_csv_dumper_276);
    mstatus_csv_dumper_277 = new("./module_status277.csv");
    module_monitor_277 = new(module_intf_277,mstatus_csv_dumper_277);
    mstatus_csv_dumper_278 = new("./module_status278.csv");
    module_monitor_278 = new(module_intf_278,mstatus_csv_dumper_278);
    mstatus_csv_dumper_279 = new("./module_status279.csv");
    module_monitor_279 = new(module_intf_279,mstatus_csv_dumper_279);
    mstatus_csv_dumper_280 = new("./module_status280.csv");
    module_monitor_280 = new(module_intf_280,mstatus_csv_dumper_280);
    mstatus_csv_dumper_281 = new("./module_status281.csv");
    module_monitor_281 = new(module_intf_281,mstatus_csv_dumper_281);
    mstatus_csv_dumper_282 = new("./module_status282.csv");
    module_monitor_282 = new(module_intf_282,mstatus_csv_dumper_282);
    mstatus_csv_dumper_283 = new("./module_status283.csv");
    module_monitor_283 = new(module_intf_283,mstatus_csv_dumper_283);
    mstatus_csv_dumper_284 = new("./module_status284.csv");
    module_monitor_284 = new(module_intf_284,mstatus_csv_dumper_284);
    mstatus_csv_dumper_285 = new("./module_status285.csv");
    module_monitor_285 = new(module_intf_285,mstatus_csv_dumper_285);
    mstatus_csv_dumper_286 = new("./module_status286.csv");
    module_monitor_286 = new(module_intf_286,mstatus_csv_dumper_286);
    mstatus_csv_dumper_287 = new("./module_status287.csv");
    module_monitor_287 = new(module_intf_287,mstatus_csv_dumper_287);
    mstatus_csv_dumper_288 = new("./module_status288.csv");
    module_monitor_288 = new(module_intf_288,mstatus_csv_dumper_288);
    mstatus_csv_dumper_289 = new("./module_status289.csv");
    module_monitor_289 = new(module_intf_289,mstatus_csv_dumper_289);
    mstatus_csv_dumper_290 = new("./module_status290.csv");
    module_monitor_290 = new(module_intf_290,mstatus_csv_dumper_290);
    mstatus_csv_dumper_291 = new("./module_status291.csv");
    module_monitor_291 = new(module_intf_291,mstatus_csv_dumper_291);
    mstatus_csv_dumper_292 = new("./module_status292.csv");
    module_monitor_292 = new(module_intf_292,mstatus_csv_dumper_292);
    mstatus_csv_dumper_293 = new("./module_status293.csv");
    module_monitor_293 = new(module_intf_293,mstatus_csv_dumper_293);
    mstatus_csv_dumper_294 = new("./module_status294.csv");
    module_monitor_294 = new(module_intf_294,mstatus_csv_dumper_294);
    mstatus_csv_dumper_295 = new("./module_status295.csv");
    module_monitor_295 = new(module_intf_295,mstatus_csv_dumper_295);
    mstatus_csv_dumper_296 = new("./module_status296.csv");
    module_monitor_296 = new(module_intf_296,mstatus_csv_dumper_296);
    mstatus_csv_dumper_297 = new("./module_status297.csv");
    module_monitor_297 = new(module_intf_297,mstatus_csv_dumper_297);
    mstatus_csv_dumper_298 = new("./module_status298.csv");
    module_monitor_298 = new(module_intf_298,mstatus_csv_dumper_298);
    mstatus_csv_dumper_299 = new("./module_status299.csv");
    module_monitor_299 = new(module_intf_299,mstatus_csv_dumper_299);
    mstatus_csv_dumper_300 = new("./module_status300.csv");
    module_monitor_300 = new(module_intf_300,mstatus_csv_dumper_300);
    mstatus_csv_dumper_301 = new("./module_status301.csv");
    module_monitor_301 = new(module_intf_301,mstatus_csv_dumper_301);
    mstatus_csv_dumper_302 = new("./module_status302.csv");
    module_monitor_302 = new(module_intf_302,mstatus_csv_dumper_302);
    mstatus_csv_dumper_303 = new("./module_status303.csv");
    module_monitor_303 = new(module_intf_303,mstatus_csv_dumper_303);
    mstatus_csv_dumper_304 = new("./module_status304.csv");
    module_monitor_304 = new(module_intf_304,mstatus_csv_dumper_304);
    mstatus_csv_dumper_305 = new("./module_status305.csv");
    module_monitor_305 = new(module_intf_305,mstatus_csv_dumper_305);
    mstatus_csv_dumper_306 = new("./module_status306.csv");
    module_monitor_306 = new(module_intf_306,mstatus_csv_dumper_306);
    mstatus_csv_dumper_307 = new("./module_status307.csv");
    module_monitor_307 = new(module_intf_307,mstatus_csv_dumper_307);
    mstatus_csv_dumper_308 = new("./module_status308.csv");
    module_monitor_308 = new(module_intf_308,mstatus_csv_dumper_308);
    mstatus_csv_dumper_309 = new("./module_status309.csv");
    module_monitor_309 = new(module_intf_309,mstatus_csv_dumper_309);
    mstatus_csv_dumper_310 = new("./module_status310.csv");
    module_monitor_310 = new(module_intf_310,mstatus_csv_dumper_310);
    mstatus_csv_dumper_311 = new("./module_status311.csv");
    module_monitor_311 = new(module_intf_311,mstatus_csv_dumper_311);
    mstatus_csv_dumper_312 = new("./module_status312.csv");
    module_monitor_312 = new(module_intf_312,mstatus_csv_dumper_312);
    mstatus_csv_dumper_313 = new("./module_status313.csv");
    module_monitor_313 = new(module_intf_313,mstatus_csv_dumper_313);
    mstatus_csv_dumper_314 = new("./module_status314.csv");
    module_monitor_314 = new(module_intf_314,mstatus_csv_dumper_314);
    mstatus_csv_dumper_315 = new("./module_status315.csv");
    module_monitor_315 = new(module_intf_315,mstatus_csv_dumper_315);
    mstatus_csv_dumper_316 = new("./module_status316.csv");
    module_monitor_316 = new(module_intf_316,mstatus_csv_dumper_316);
    mstatus_csv_dumper_317 = new("./module_status317.csv");
    module_monitor_317 = new(module_intf_317,mstatus_csv_dumper_317);
    mstatus_csv_dumper_318 = new("./module_status318.csv");
    module_monitor_318 = new(module_intf_318,mstatus_csv_dumper_318);
    mstatus_csv_dumper_319 = new("./module_status319.csv");
    module_monitor_319 = new(module_intf_319,mstatus_csv_dumper_319);
    mstatus_csv_dumper_320 = new("./module_status320.csv");
    module_monitor_320 = new(module_intf_320,mstatus_csv_dumper_320);
    mstatus_csv_dumper_321 = new("./module_status321.csv");
    module_monitor_321 = new(module_intf_321,mstatus_csv_dumper_321);
    mstatus_csv_dumper_322 = new("./module_status322.csv");
    module_monitor_322 = new(module_intf_322,mstatus_csv_dumper_322);
    mstatus_csv_dumper_323 = new("./module_status323.csv");
    module_monitor_323 = new(module_intf_323,mstatus_csv_dumper_323);
    mstatus_csv_dumper_324 = new("./module_status324.csv");
    module_monitor_324 = new(module_intf_324,mstatus_csv_dumper_324);
    mstatus_csv_dumper_325 = new("./module_status325.csv");
    module_monitor_325 = new(module_intf_325,mstatus_csv_dumper_325);
    mstatus_csv_dumper_326 = new("./module_status326.csv");
    module_monitor_326 = new(module_intf_326,mstatus_csv_dumper_326);
    mstatus_csv_dumper_327 = new("./module_status327.csv");
    module_monitor_327 = new(module_intf_327,mstatus_csv_dumper_327);
    mstatus_csv_dumper_328 = new("./module_status328.csv");
    module_monitor_328 = new(module_intf_328,mstatus_csv_dumper_328);
    mstatus_csv_dumper_329 = new("./module_status329.csv");
    module_monitor_329 = new(module_intf_329,mstatus_csv_dumper_329);
    mstatus_csv_dumper_330 = new("./module_status330.csv");
    module_monitor_330 = new(module_intf_330,mstatus_csv_dumper_330);
    mstatus_csv_dumper_331 = new("./module_status331.csv");
    module_monitor_331 = new(module_intf_331,mstatus_csv_dumper_331);
    mstatus_csv_dumper_332 = new("./module_status332.csv");
    module_monitor_332 = new(module_intf_332,mstatus_csv_dumper_332);
    mstatus_csv_dumper_333 = new("./module_status333.csv");
    module_monitor_333 = new(module_intf_333,mstatus_csv_dumper_333);
    mstatus_csv_dumper_334 = new("./module_status334.csv");
    module_monitor_334 = new(module_intf_334,mstatus_csv_dumper_334);
    mstatus_csv_dumper_335 = new("./module_status335.csv");
    module_monitor_335 = new(module_intf_335,mstatus_csv_dumper_335);
    mstatus_csv_dumper_336 = new("./module_status336.csv");
    module_monitor_336 = new(module_intf_336,mstatus_csv_dumper_336);
    mstatus_csv_dumper_337 = new("./module_status337.csv");
    module_monitor_337 = new(module_intf_337,mstatus_csv_dumper_337);
    mstatus_csv_dumper_338 = new("./module_status338.csv");
    module_monitor_338 = new(module_intf_338,mstatus_csv_dumper_338);
    mstatus_csv_dumper_339 = new("./module_status339.csv");
    module_monitor_339 = new(module_intf_339,mstatus_csv_dumper_339);
    mstatus_csv_dumper_340 = new("./module_status340.csv");
    module_monitor_340 = new(module_intf_340,mstatus_csv_dumper_340);
    mstatus_csv_dumper_341 = new("./module_status341.csv");
    module_monitor_341 = new(module_intf_341,mstatus_csv_dumper_341);
    mstatus_csv_dumper_342 = new("./module_status342.csv");
    module_monitor_342 = new(module_intf_342,mstatus_csv_dumper_342);
    mstatus_csv_dumper_343 = new("./module_status343.csv");
    module_monitor_343 = new(module_intf_343,mstatus_csv_dumper_343);
    mstatus_csv_dumper_344 = new("./module_status344.csv");
    module_monitor_344 = new(module_intf_344,mstatus_csv_dumper_344);
    mstatus_csv_dumper_345 = new("./module_status345.csv");
    module_monitor_345 = new(module_intf_345,mstatus_csv_dumper_345);
    mstatus_csv_dumper_346 = new("./module_status346.csv");
    module_monitor_346 = new(module_intf_346,mstatus_csv_dumper_346);
    mstatus_csv_dumper_347 = new("./module_status347.csv");
    module_monitor_347 = new(module_intf_347,mstatus_csv_dumper_347);
    mstatus_csv_dumper_348 = new("./module_status348.csv");
    module_monitor_348 = new(module_intf_348,mstatus_csv_dumper_348);
    mstatus_csv_dumper_349 = new("./module_status349.csv");
    module_monitor_349 = new(module_intf_349,mstatus_csv_dumper_349);
    mstatus_csv_dumper_350 = new("./module_status350.csv");
    module_monitor_350 = new(module_intf_350,mstatus_csv_dumper_350);
    mstatus_csv_dumper_351 = new("./module_status351.csv");
    module_monitor_351 = new(module_intf_351,mstatus_csv_dumper_351);
    mstatus_csv_dumper_352 = new("./module_status352.csv");
    module_monitor_352 = new(module_intf_352,mstatus_csv_dumper_352);
    mstatus_csv_dumper_353 = new("./module_status353.csv");
    module_monitor_353 = new(module_intf_353,mstatus_csv_dumper_353);
    mstatus_csv_dumper_354 = new("./module_status354.csv");
    module_monitor_354 = new(module_intf_354,mstatus_csv_dumper_354);
    mstatus_csv_dumper_355 = new("./module_status355.csv");
    module_monitor_355 = new(module_intf_355,mstatus_csv_dumper_355);
    mstatus_csv_dumper_356 = new("./module_status356.csv");
    module_monitor_356 = new(module_intf_356,mstatus_csv_dumper_356);
    mstatus_csv_dumper_357 = new("./module_status357.csv");
    module_monitor_357 = new(module_intf_357,mstatus_csv_dumper_357);
    mstatus_csv_dumper_358 = new("./module_status358.csv");
    module_monitor_358 = new(module_intf_358,mstatus_csv_dumper_358);
    mstatus_csv_dumper_359 = new("./module_status359.csv");
    module_monitor_359 = new(module_intf_359,mstatus_csv_dumper_359);
    mstatus_csv_dumper_360 = new("./module_status360.csv");
    module_monitor_360 = new(module_intf_360,mstatus_csv_dumper_360);
    mstatus_csv_dumper_361 = new("./module_status361.csv");
    module_monitor_361 = new(module_intf_361,mstatus_csv_dumper_361);
    mstatus_csv_dumper_362 = new("./module_status362.csv");
    module_monitor_362 = new(module_intf_362,mstatus_csv_dumper_362);
    mstatus_csv_dumper_363 = new("./module_status363.csv");
    module_monitor_363 = new(module_intf_363,mstatus_csv_dumper_363);
    mstatus_csv_dumper_364 = new("./module_status364.csv");
    module_monitor_364 = new(module_intf_364,mstatus_csv_dumper_364);
    mstatus_csv_dumper_365 = new("./module_status365.csv");
    module_monitor_365 = new(module_intf_365,mstatus_csv_dumper_365);
    mstatus_csv_dumper_366 = new("./module_status366.csv");
    module_monitor_366 = new(module_intf_366,mstatus_csv_dumper_366);
    mstatus_csv_dumper_367 = new("./module_status367.csv");
    module_monitor_367 = new(module_intf_367,mstatus_csv_dumper_367);
    mstatus_csv_dumper_368 = new("./module_status368.csv");
    module_monitor_368 = new(module_intf_368,mstatus_csv_dumper_368);
    mstatus_csv_dumper_369 = new("./module_status369.csv");
    module_monitor_369 = new(module_intf_369,mstatus_csv_dumper_369);
    mstatus_csv_dumper_370 = new("./module_status370.csv");
    module_monitor_370 = new(module_intf_370,mstatus_csv_dumper_370);
    mstatus_csv_dumper_371 = new("./module_status371.csv");
    module_monitor_371 = new(module_intf_371,mstatus_csv_dumper_371);
    mstatus_csv_dumper_372 = new("./module_status372.csv");
    module_monitor_372 = new(module_intf_372,mstatus_csv_dumper_372);
    mstatus_csv_dumper_373 = new("./module_status373.csv");
    module_monitor_373 = new(module_intf_373,mstatus_csv_dumper_373);
    mstatus_csv_dumper_374 = new("./module_status374.csv");
    module_monitor_374 = new(module_intf_374,mstatus_csv_dumper_374);
    mstatus_csv_dumper_375 = new("./module_status375.csv");
    module_monitor_375 = new(module_intf_375,mstatus_csv_dumper_375);
    mstatus_csv_dumper_376 = new("./module_status376.csv");
    module_monitor_376 = new(module_intf_376,mstatus_csv_dumper_376);
    mstatus_csv_dumper_377 = new("./module_status377.csv");
    module_monitor_377 = new(module_intf_377,mstatus_csv_dumper_377);
    mstatus_csv_dumper_378 = new("./module_status378.csv");
    module_monitor_378 = new(module_intf_378,mstatus_csv_dumper_378);
    mstatus_csv_dumper_379 = new("./module_status379.csv");
    module_monitor_379 = new(module_intf_379,mstatus_csv_dumper_379);
    mstatus_csv_dumper_380 = new("./module_status380.csv");
    module_monitor_380 = new(module_intf_380,mstatus_csv_dumper_380);
    mstatus_csv_dumper_381 = new("./module_status381.csv");
    module_monitor_381 = new(module_intf_381,mstatus_csv_dumper_381);
    mstatus_csv_dumper_382 = new("./module_status382.csv");
    module_monitor_382 = new(module_intf_382,mstatus_csv_dumper_382);
    mstatus_csv_dumper_383 = new("./module_status383.csv");
    module_monitor_383 = new(module_intf_383,mstatus_csv_dumper_383);
    mstatus_csv_dumper_384 = new("./module_status384.csv");
    module_monitor_384 = new(module_intf_384,mstatus_csv_dumper_384);
    mstatus_csv_dumper_385 = new("./module_status385.csv");
    module_monitor_385 = new(module_intf_385,mstatus_csv_dumper_385);
    mstatus_csv_dumper_386 = new("./module_status386.csv");
    module_monitor_386 = new(module_intf_386,mstatus_csv_dumper_386);
    mstatus_csv_dumper_387 = new("./module_status387.csv");
    module_monitor_387 = new(module_intf_387,mstatus_csv_dumper_387);
    mstatus_csv_dumper_388 = new("./module_status388.csv");
    module_monitor_388 = new(module_intf_388,mstatus_csv_dumper_388);
    mstatus_csv_dumper_389 = new("./module_status389.csv");
    module_monitor_389 = new(module_intf_389,mstatus_csv_dumper_389);
    mstatus_csv_dumper_390 = new("./module_status390.csv");
    module_monitor_390 = new(module_intf_390,mstatus_csv_dumper_390);
    mstatus_csv_dumper_391 = new("./module_status391.csv");
    module_monitor_391 = new(module_intf_391,mstatus_csv_dumper_391);
    mstatus_csv_dumper_392 = new("./module_status392.csv");
    module_monitor_392 = new(module_intf_392,mstatus_csv_dumper_392);
    mstatus_csv_dumper_393 = new("./module_status393.csv");
    module_monitor_393 = new(module_intf_393,mstatus_csv_dumper_393);
    mstatus_csv_dumper_394 = new("./module_status394.csv");
    module_monitor_394 = new(module_intf_394,mstatus_csv_dumper_394);
    mstatus_csv_dumper_395 = new("./module_status395.csv");
    module_monitor_395 = new(module_intf_395,mstatus_csv_dumper_395);
    mstatus_csv_dumper_396 = new("./module_status396.csv");
    module_monitor_396 = new(module_intf_396,mstatus_csv_dumper_396);
    mstatus_csv_dumper_397 = new("./module_status397.csv");
    module_monitor_397 = new(module_intf_397,mstatus_csv_dumper_397);
    mstatus_csv_dumper_398 = new("./module_status398.csv");
    module_monitor_398 = new(module_intf_398,mstatus_csv_dumper_398);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    sample_manager_inst.add_one_monitor(module_monitor_58);
    sample_manager_inst.add_one_monitor(module_monitor_59);
    sample_manager_inst.add_one_monitor(module_monitor_60);
    sample_manager_inst.add_one_monitor(module_monitor_61);
    sample_manager_inst.add_one_monitor(module_monitor_62);
    sample_manager_inst.add_one_monitor(module_monitor_63);
    sample_manager_inst.add_one_monitor(module_monitor_64);
    sample_manager_inst.add_one_monitor(module_monitor_65);
    sample_manager_inst.add_one_monitor(module_monitor_66);
    sample_manager_inst.add_one_monitor(module_monitor_67);
    sample_manager_inst.add_one_monitor(module_monitor_68);
    sample_manager_inst.add_one_monitor(module_monitor_69);
    sample_manager_inst.add_one_monitor(module_monitor_70);
    sample_manager_inst.add_one_monitor(module_monitor_71);
    sample_manager_inst.add_one_monitor(module_monitor_72);
    sample_manager_inst.add_one_monitor(module_monitor_73);
    sample_manager_inst.add_one_monitor(module_monitor_74);
    sample_manager_inst.add_one_monitor(module_monitor_75);
    sample_manager_inst.add_one_monitor(module_monitor_76);
    sample_manager_inst.add_one_monitor(module_monitor_77);
    sample_manager_inst.add_one_monitor(module_monitor_78);
    sample_manager_inst.add_one_monitor(module_monitor_79);
    sample_manager_inst.add_one_monitor(module_monitor_80);
    sample_manager_inst.add_one_monitor(module_monitor_81);
    sample_manager_inst.add_one_monitor(module_monitor_82);
    sample_manager_inst.add_one_monitor(module_monitor_83);
    sample_manager_inst.add_one_monitor(module_monitor_84);
    sample_manager_inst.add_one_monitor(module_monitor_85);
    sample_manager_inst.add_one_monitor(module_monitor_86);
    sample_manager_inst.add_one_monitor(module_monitor_87);
    sample_manager_inst.add_one_monitor(module_monitor_88);
    sample_manager_inst.add_one_monitor(module_monitor_89);
    sample_manager_inst.add_one_monitor(module_monitor_90);
    sample_manager_inst.add_one_monitor(module_monitor_91);
    sample_manager_inst.add_one_monitor(module_monitor_92);
    sample_manager_inst.add_one_monitor(module_monitor_93);
    sample_manager_inst.add_one_monitor(module_monitor_94);
    sample_manager_inst.add_one_monitor(module_monitor_95);
    sample_manager_inst.add_one_monitor(module_monitor_96);
    sample_manager_inst.add_one_monitor(module_monitor_97);
    sample_manager_inst.add_one_monitor(module_monitor_98);
    sample_manager_inst.add_one_monitor(module_monitor_99);
    sample_manager_inst.add_one_monitor(module_monitor_100);
    sample_manager_inst.add_one_monitor(module_monitor_101);
    sample_manager_inst.add_one_monitor(module_monitor_102);
    sample_manager_inst.add_one_monitor(module_monitor_103);
    sample_manager_inst.add_one_monitor(module_monitor_104);
    sample_manager_inst.add_one_monitor(module_monitor_105);
    sample_manager_inst.add_one_monitor(module_monitor_106);
    sample_manager_inst.add_one_monitor(module_monitor_107);
    sample_manager_inst.add_one_monitor(module_monitor_108);
    sample_manager_inst.add_one_monitor(module_monitor_109);
    sample_manager_inst.add_one_monitor(module_monitor_110);
    sample_manager_inst.add_one_monitor(module_monitor_111);
    sample_manager_inst.add_one_monitor(module_monitor_112);
    sample_manager_inst.add_one_monitor(module_monitor_113);
    sample_manager_inst.add_one_monitor(module_monitor_114);
    sample_manager_inst.add_one_monitor(module_monitor_115);
    sample_manager_inst.add_one_monitor(module_monitor_116);
    sample_manager_inst.add_one_monitor(module_monitor_117);
    sample_manager_inst.add_one_monitor(module_monitor_118);
    sample_manager_inst.add_one_monitor(module_monitor_119);
    sample_manager_inst.add_one_monitor(module_monitor_120);
    sample_manager_inst.add_one_monitor(module_monitor_121);
    sample_manager_inst.add_one_monitor(module_monitor_122);
    sample_manager_inst.add_one_monitor(module_monitor_123);
    sample_manager_inst.add_one_monitor(module_monitor_124);
    sample_manager_inst.add_one_monitor(module_monitor_125);
    sample_manager_inst.add_one_monitor(module_monitor_126);
    sample_manager_inst.add_one_monitor(module_monitor_127);
    sample_manager_inst.add_one_monitor(module_monitor_128);
    sample_manager_inst.add_one_monitor(module_monitor_129);
    sample_manager_inst.add_one_monitor(module_monitor_130);
    sample_manager_inst.add_one_monitor(module_monitor_131);
    sample_manager_inst.add_one_monitor(module_monitor_132);
    sample_manager_inst.add_one_monitor(module_monitor_133);
    sample_manager_inst.add_one_monitor(module_monitor_134);
    sample_manager_inst.add_one_monitor(module_monitor_135);
    sample_manager_inst.add_one_monitor(module_monitor_136);
    sample_manager_inst.add_one_monitor(module_monitor_137);
    sample_manager_inst.add_one_monitor(module_monitor_138);
    sample_manager_inst.add_one_monitor(module_monitor_139);
    sample_manager_inst.add_one_monitor(module_monitor_140);
    sample_manager_inst.add_one_monitor(module_monitor_141);
    sample_manager_inst.add_one_monitor(module_monitor_142);
    sample_manager_inst.add_one_monitor(module_monitor_143);
    sample_manager_inst.add_one_monitor(module_monitor_144);
    sample_manager_inst.add_one_monitor(module_monitor_145);
    sample_manager_inst.add_one_monitor(module_monitor_146);
    sample_manager_inst.add_one_monitor(module_monitor_147);
    sample_manager_inst.add_one_monitor(module_monitor_148);
    sample_manager_inst.add_one_monitor(module_monitor_149);
    sample_manager_inst.add_one_monitor(module_monitor_150);
    sample_manager_inst.add_one_monitor(module_monitor_151);
    sample_manager_inst.add_one_monitor(module_monitor_152);
    sample_manager_inst.add_one_monitor(module_monitor_153);
    sample_manager_inst.add_one_monitor(module_monitor_154);
    sample_manager_inst.add_one_monitor(module_monitor_155);
    sample_manager_inst.add_one_monitor(module_monitor_156);
    sample_manager_inst.add_one_monitor(module_monitor_157);
    sample_manager_inst.add_one_monitor(module_monitor_158);
    sample_manager_inst.add_one_monitor(module_monitor_159);
    sample_manager_inst.add_one_monitor(module_monitor_160);
    sample_manager_inst.add_one_monitor(module_monitor_161);
    sample_manager_inst.add_one_monitor(module_monitor_162);
    sample_manager_inst.add_one_monitor(module_monitor_163);
    sample_manager_inst.add_one_monitor(module_monitor_164);
    sample_manager_inst.add_one_monitor(module_monitor_165);
    sample_manager_inst.add_one_monitor(module_monitor_166);
    sample_manager_inst.add_one_monitor(module_monitor_167);
    sample_manager_inst.add_one_monitor(module_monitor_168);
    sample_manager_inst.add_one_monitor(module_monitor_169);
    sample_manager_inst.add_one_monitor(module_monitor_170);
    sample_manager_inst.add_one_monitor(module_monitor_171);
    sample_manager_inst.add_one_monitor(module_monitor_172);
    sample_manager_inst.add_one_monitor(module_monitor_173);
    sample_manager_inst.add_one_monitor(module_monitor_174);
    sample_manager_inst.add_one_monitor(module_monitor_175);
    sample_manager_inst.add_one_monitor(module_monitor_176);
    sample_manager_inst.add_one_monitor(module_monitor_177);
    sample_manager_inst.add_one_monitor(module_monitor_178);
    sample_manager_inst.add_one_monitor(module_monitor_179);
    sample_manager_inst.add_one_monitor(module_monitor_180);
    sample_manager_inst.add_one_monitor(module_monitor_181);
    sample_manager_inst.add_one_monitor(module_monitor_182);
    sample_manager_inst.add_one_monitor(module_monitor_183);
    sample_manager_inst.add_one_monitor(module_monitor_184);
    sample_manager_inst.add_one_monitor(module_monitor_185);
    sample_manager_inst.add_one_monitor(module_monitor_186);
    sample_manager_inst.add_one_monitor(module_monitor_187);
    sample_manager_inst.add_one_monitor(module_monitor_188);
    sample_manager_inst.add_one_monitor(module_monitor_189);
    sample_manager_inst.add_one_monitor(module_monitor_190);
    sample_manager_inst.add_one_monitor(module_monitor_191);
    sample_manager_inst.add_one_monitor(module_monitor_192);
    sample_manager_inst.add_one_monitor(module_monitor_193);
    sample_manager_inst.add_one_monitor(module_monitor_194);
    sample_manager_inst.add_one_monitor(module_monitor_195);
    sample_manager_inst.add_one_monitor(module_monitor_196);
    sample_manager_inst.add_one_monitor(module_monitor_197);
    sample_manager_inst.add_one_monitor(module_monitor_198);
    sample_manager_inst.add_one_monitor(module_monitor_199);
    sample_manager_inst.add_one_monitor(module_monitor_200);
    sample_manager_inst.add_one_monitor(module_monitor_201);
    sample_manager_inst.add_one_monitor(module_monitor_202);
    sample_manager_inst.add_one_monitor(module_monitor_203);
    sample_manager_inst.add_one_monitor(module_monitor_204);
    sample_manager_inst.add_one_monitor(module_monitor_205);
    sample_manager_inst.add_one_monitor(module_monitor_206);
    sample_manager_inst.add_one_monitor(module_monitor_207);
    sample_manager_inst.add_one_monitor(module_monitor_208);
    sample_manager_inst.add_one_monitor(module_monitor_209);
    sample_manager_inst.add_one_monitor(module_monitor_210);
    sample_manager_inst.add_one_monitor(module_monitor_211);
    sample_manager_inst.add_one_monitor(module_monitor_212);
    sample_manager_inst.add_one_monitor(module_monitor_213);
    sample_manager_inst.add_one_monitor(module_monitor_214);
    sample_manager_inst.add_one_monitor(module_monitor_215);
    sample_manager_inst.add_one_monitor(module_monitor_216);
    sample_manager_inst.add_one_monitor(module_monitor_217);
    sample_manager_inst.add_one_monitor(module_monitor_218);
    sample_manager_inst.add_one_monitor(module_monitor_219);
    sample_manager_inst.add_one_monitor(module_monitor_220);
    sample_manager_inst.add_one_monitor(module_monitor_221);
    sample_manager_inst.add_one_monitor(module_monitor_222);
    sample_manager_inst.add_one_monitor(module_monitor_223);
    sample_manager_inst.add_one_monitor(module_monitor_224);
    sample_manager_inst.add_one_monitor(module_monitor_225);
    sample_manager_inst.add_one_monitor(module_monitor_226);
    sample_manager_inst.add_one_monitor(module_monitor_227);
    sample_manager_inst.add_one_monitor(module_monitor_228);
    sample_manager_inst.add_one_monitor(module_monitor_229);
    sample_manager_inst.add_one_monitor(module_monitor_230);
    sample_manager_inst.add_one_monitor(module_monitor_231);
    sample_manager_inst.add_one_monitor(module_monitor_232);
    sample_manager_inst.add_one_monitor(module_monitor_233);
    sample_manager_inst.add_one_monitor(module_monitor_234);
    sample_manager_inst.add_one_monitor(module_monitor_235);
    sample_manager_inst.add_one_monitor(module_monitor_236);
    sample_manager_inst.add_one_monitor(module_monitor_237);
    sample_manager_inst.add_one_monitor(module_monitor_238);
    sample_manager_inst.add_one_monitor(module_monitor_239);
    sample_manager_inst.add_one_monitor(module_monitor_240);
    sample_manager_inst.add_one_monitor(module_monitor_241);
    sample_manager_inst.add_one_monitor(module_monitor_242);
    sample_manager_inst.add_one_monitor(module_monitor_243);
    sample_manager_inst.add_one_monitor(module_monitor_244);
    sample_manager_inst.add_one_monitor(module_monitor_245);
    sample_manager_inst.add_one_monitor(module_monitor_246);
    sample_manager_inst.add_one_monitor(module_monitor_247);
    sample_manager_inst.add_one_monitor(module_monitor_248);
    sample_manager_inst.add_one_monitor(module_monitor_249);
    sample_manager_inst.add_one_monitor(module_monitor_250);
    sample_manager_inst.add_one_monitor(module_monitor_251);
    sample_manager_inst.add_one_monitor(module_monitor_252);
    sample_manager_inst.add_one_monitor(module_monitor_253);
    sample_manager_inst.add_one_monitor(module_monitor_254);
    sample_manager_inst.add_one_monitor(module_monitor_255);
    sample_manager_inst.add_one_monitor(module_monitor_256);
    sample_manager_inst.add_one_monitor(module_monitor_257);
    sample_manager_inst.add_one_monitor(module_monitor_258);
    sample_manager_inst.add_one_monitor(module_monitor_259);
    sample_manager_inst.add_one_monitor(module_monitor_260);
    sample_manager_inst.add_one_monitor(module_monitor_261);
    sample_manager_inst.add_one_monitor(module_monitor_262);
    sample_manager_inst.add_one_monitor(module_monitor_263);
    sample_manager_inst.add_one_monitor(module_monitor_264);
    sample_manager_inst.add_one_monitor(module_monitor_265);
    sample_manager_inst.add_one_monitor(module_monitor_266);
    sample_manager_inst.add_one_monitor(module_monitor_267);
    sample_manager_inst.add_one_monitor(module_monitor_268);
    sample_manager_inst.add_one_monitor(module_monitor_269);
    sample_manager_inst.add_one_monitor(module_monitor_270);
    sample_manager_inst.add_one_monitor(module_monitor_271);
    sample_manager_inst.add_one_monitor(module_monitor_272);
    sample_manager_inst.add_one_monitor(module_monitor_273);
    sample_manager_inst.add_one_monitor(module_monitor_274);
    sample_manager_inst.add_one_monitor(module_monitor_275);
    sample_manager_inst.add_one_monitor(module_monitor_276);
    sample_manager_inst.add_one_monitor(module_monitor_277);
    sample_manager_inst.add_one_monitor(module_monitor_278);
    sample_manager_inst.add_one_monitor(module_monitor_279);
    sample_manager_inst.add_one_monitor(module_monitor_280);
    sample_manager_inst.add_one_monitor(module_monitor_281);
    sample_manager_inst.add_one_monitor(module_monitor_282);
    sample_manager_inst.add_one_monitor(module_monitor_283);
    sample_manager_inst.add_one_monitor(module_monitor_284);
    sample_manager_inst.add_one_monitor(module_monitor_285);
    sample_manager_inst.add_one_monitor(module_monitor_286);
    sample_manager_inst.add_one_monitor(module_monitor_287);
    sample_manager_inst.add_one_monitor(module_monitor_288);
    sample_manager_inst.add_one_monitor(module_monitor_289);
    sample_manager_inst.add_one_monitor(module_monitor_290);
    sample_manager_inst.add_one_monitor(module_monitor_291);
    sample_manager_inst.add_one_monitor(module_monitor_292);
    sample_manager_inst.add_one_monitor(module_monitor_293);
    sample_manager_inst.add_one_monitor(module_monitor_294);
    sample_manager_inst.add_one_monitor(module_monitor_295);
    sample_manager_inst.add_one_monitor(module_monitor_296);
    sample_manager_inst.add_one_monitor(module_monitor_297);
    sample_manager_inst.add_one_monitor(module_monitor_298);
    sample_manager_inst.add_one_monitor(module_monitor_299);
    sample_manager_inst.add_one_monitor(module_monitor_300);
    sample_manager_inst.add_one_monitor(module_monitor_301);
    sample_manager_inst.add_one_monitor(module_monitor_302);
    sample_manager_inst.add_one_monitor(module_monitor_303);
    sample_manager_inst.add_one_monitor(module_monitor_304);
    sample_manager_inst.add_one_monitor(module_monitor_305);
    sample_manager_inst.add_one_monitor(module_monitor_306);
    sample_manager_inst.add_one_monitor(module_monitor_307);
    sample_manager_inst.add_one_monitor(module_monitor_308);
    sample_manager_inst.add_one_monitor(module_monitor_309);
    sample_manager_inst.add_one_monitor(module_monitor_310);
    sample_manager_inst.add_one_monitor(module_monitor_311);
    sample_manager_inst.add_one_monitor(module_monitor_312);
    sample_manager_inst.add_one_monitor(module_monitor_313);
    sample_manager_inst.add_one_monitor(module_monitor_314);
    sample_manager_inst.add_one_monitor(module_monitor_315);
    sample_manager_inst.add_one_monitor(module_monitor_316);
    sample_manager_inst.add_one_monitor(module_monitor_317);
    sample_manager_inst.add_one_monitor(module_monitor_318);
    sample_manager_inst.add_one_monitor(module_monitor_319);
    sample_manager_inst.add_one_monitor(module_monitor_320);
    sample_manager_inst.add_one_monitor(module_monitor_321);
    sample_manager_inst.add_one_monitor(module_monitor_322);
    sample_manager_inst.add_one_monitor(module_monitor_323);
    sample_manager_inst.add_one_monitor(module_monitor_324);
    sample_manager_inst.add_one_monitor(module_monitor_325);
    sample_manager_inst.add_one_monitor(module_monitor_326);
    sample_manager_inst.add_one_monitor(module_monitor_327);
    sample_manager_inst.add_one_monitor(module_monitor_328);
    sample_manager_inst.add_one_monitor(module_monitor_329);
    sample_manager_inst.add_one_monitor(module_monitor_330);
    sample_manager_inst.add_one_monitor(module_monitor_331);
    sample_manager_inst.add_one_monitor(module_monitor_332);
    sample_manager_inst.add_one_monitor(module_monitor_333);
    sample_manager_inst.add_one_monitor(module_monitor_334);
    sample_manager_inst.add_one_monitor(module_monitor_335);
    sample_manager_inst.add_one_monitor(module_monitor_336);
    sample_manager_inst.add_one_monitor(module_monitor_337);
    sample_manager_inst.add_one_monitor(module_monitor_338);
    sample_manager_inst.add_one_monitor(module_monitor_339);
    sample_manager_inst.add_one_monitor(module_monitor_340);
    sample_manager_inst.add_one_monitor(module_monitor_341);
    sample_manager_inst.add_one_monitor(module_monitor_342);
    sample_manager_inst.add_one_monitor(module_monitor_343);
    sample_manager_inst.add_one_monitor(module_monitor_344);
    sample_manager_inst.add_one_monitor(module_monitor_345);
    sample_manager_inst.add_one_monitor(module_monitor_346);
    sample_manager_inst.add_one_monitor(module_monitor_347);
    sample_manager_inst.add_one_monitor(module_monitor_348);
    sample_manager_inst.add_one_monitor(module_monitor_349);
    sample_manager_inst.add_one_monitor(module_monitor_350);
    sample_manager_inst.add_one_monitor(module_monitor_351);
    sample_manager_inst.add_one_monitor(module_monitor_352);
    sample_manager_inst.add_one_monitor(module_monitor_353);
    sample_manager_inst.add_one_monitor(module_monitor_354);
    sample_manager_inst.add_one_monitor(module_monitor_355);
    sample_manager_inst.add_one_monitor(module_monitor_356);
    sample_manager_inst.add_one_monitor(module_monitor_357);
    sample_manager_inst.add_one_monitor(module_monitor_358);
    sample_manager_inst.add_one_monitor(module_monitor_359);
    sample_manager_inst.add_one_monitor(module_monitor_360);
    sample_manager_inst.add_one_monitor(module_monitor_361);
    sample_manager_inst.add_one_monitor(module_monitor_362);
    sample_manager_inst.add_one_monitor(module_monitor_363);
    sample_manager_inst.add_one_monitor(module_monitor_364);
    sample_manager_inst.add_one_monitor(module_monitor_365);
    sample_manager_inst.add_one_monitor(module_monitor_366);
    sample_manager_inst.add_one_monitor(module_monitor_367);
    sample_manager_inst.add_one_monitor(module_monitor_368);
    sample_manager_inst.add_one_monitor(module_monitor_369);
    sample_manager_inst.add_one_monitor(module_monitor_370);
    sample_manager_inst.add_one_monitor(module_monitor_371);
    sample_manager_inst.add_one_monitor(module_monitor_372);
    sample_manager_inst.add_one_monitor(module_monitor_373);
    sample_manager_inst.add_one_monitor(module_monitor_374);
    sample_manager_inst.add_one_monitor(module_monitor_375);
    sample_manager_inst.add_one_monitor(module_monitor_376);
    sample_manager_inst.add_one_monitor(module_monitor_377);
    sample_manager_inst.add_one_monitor(module_monitor_378);
    sample_manager_inst.add_one_monitor(module_monitor_379);
    sample_manager_inst.add_one_monitor(module_monitor_380);
    sample_manager_inst.add_one_monitor(module_monitor_381);
    sample_manager_inst.add_one_monitor(module_monitor_382);
    sample_manager_inst.add_one_monitor(module_monitor_383);
    sample_manager_inst.add_one_monitor(module_monitor_384);
    sample_manager_inst.add_one_monitor(module_monitor_385);
    sample_manager_inst.add_one_monitor(module_monitor_386);
    sample_manager_inst.add_one_monitor(module_monitor_387);
    sample_manager_inst.add_one_monitor(module_monitor_388);
    sample_manager_inst.add_one_monitor(module_monitor_389);
    sample_manager_inst.add_one_monitor(module_monitor_390);
    sample_manager_inst.add_one_monitor(module_monitor_391);
    sample_manager_inst.add_one_monitor(module_monitor_392);
    sample_manager_inst.add_one_monitor(module_monitor_393);
    sample_manager_inst.add_one_monitor(module_monitor_394);
    sample_manager_inst.add_one_monitor(module_monitor_395);
    sample_manager_inst.add_one_monitor(module_monitor_396);
    sample_manager_inst.add_one_monitor(module_monitor_397);
    sample_manager_inst.add_one_monitor(module_monitor_398);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
