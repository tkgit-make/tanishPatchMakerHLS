
`include "sample_manager.sv"
`include "csv_file_dump.sv"
`include "df_fifo_monitor.sv"
`include "df_process_monitor.sv"
`include "nodf_module_monitor.sv"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_MPSQ.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_MPSQ.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_MPSQ.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_add_patch9_fu_433.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_add_patch9_fu_433.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_add_patch9_fu_433.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = 1'b0;
    assign module_intf_17.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_makePatch_alignedToLine_fu_494.grp_add_patch9_fu_433.grp_encodeCoordinates_fu_494.ap_ready;
    assign module_intf_17.ap_done = 1'b0;
    assign module_intf_17.ap_continue = 1'b0;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_getShadows_fu_517.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_getShadows_fu_517.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_getShadows_fu_517.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_getShadows_fu_517.grp_straightLineProjectorFromLayerIJtoK_fu_245.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_getShadows_fu_517.grp_straightLineProjectorFromLayerIJtoK_fu_245.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_getShadows_fu_517.grp_straightLineProjectorFromLayerIJtoK_fu_245.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_delete_patch_fu_533.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_delete_patch_fu_533.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makeThirdPatch_fu_481.grp_delete_patch_fu_533.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_add_patch9_fu_433.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_add_patch9_fu_433.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_add_patch9_fu_433.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = 1'b0;
    assign module_intf_34.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_makePatch_alignedToLine_fu_649.grp_add_patch9_fu_433.grp_encodeCoordinates_fu_494.ap_ready;
    assign module_intf_34.ap_done = 1'b0;
    assign module_intf_34.ap_continue = 1'b0;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_delete_patch_fu_672.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_delete_patch_fu_672.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_delete_patch_fu_672.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_get_index_from_z_fu_698.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_get_index_from_z_fu_698.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_get_index_from_z_fu_698.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_areWedgeSuperPointsEqual_fu_712.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_areWedgeSuperPointsEqual_fu_712.ap_ready;
    assign module_intf_37.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_solveComplmentaryPatch_fu_508.grp_areWedgeSuperPointsEqual_fu_712.ap_done;
    assign module_intf_37.ap_continue = 1'b1;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_ready;
    assign module_intf_41.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_202.ap_done;
    assign module_intf_41.ap_continue = 1'b1;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_215.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_228.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_ready;
    assign module_intf_44.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_getParallelograms_fu_239.grp_straightLineProjectorFromLayerIJtoK_fu_241.ap_done;
    assign module_intf_44.ap_continue = 1'b1;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_wedgePatch_init_fu_404.grp_get_acceptanceCorners_fu_249.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findLRBounds_fu_282.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_ready;
    assign module_intf_48.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_makeSuperPoint_alignedToLine11_fu_414.grp_mSP_findStartIndex_fu_292.ap_done;
    assign module_intf_48.ap_continue = 1'b1;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_add_patch9_fu_433.ap_start;
    assign module_intf_49.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_add_patch9_fu_433.ap_ready;
    assign module_intf_49.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_add_patch9_fu_433.ap_done;
    assign module_intf_49.ap_continue = 1'b1;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = 1'b0;
    assign module_intf_50.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_makePatch_alignedToLine_fu_541.grp_add_patch9_fu_433.grp_encodeCoordinates_fu_494.ap_ready;
    assign module_intf_50.ap_done = 1'b0;
    assign module_intf_50.ap_continue = 1'b0;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_straightLineProjectorFromLayerIJtoK_fu_568.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_straightLineProjectorFromLayerIJtoK_fu_568.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_straightLineProjectorFromLayerIJtoK_fu_568.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_getSolveNextPatchPairWhileCondition_fu_582.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_getSolveNextPatchPairWhileCondition_fu_582.ap_ready;
    assign module_intf_52.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_getSolveNextPatchPairWhileCondition_fu_582.ap_done;
    assign module_intf_52.ap_continue = 1'b1;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_areWedgeSuperPointsEqual_fu_600.ap_start;
    assign module_intf_53.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_areWedgeSuperPointsEqual_fu_600.ap_ready;
    assign module_intf_53.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_areWedgeSuperPointsEqual_fu_600.ap_done;
    assign module_intf_53.ap_continue = 1'b1;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_straightLineProjectorFromLayerIJtoK_fu_1464.ap_start;
    assign module_intf_54.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_straightLineProjectorFromLayerIJtoK_fu_1464.ap_ready;
    assign module_intf_54.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_solveNextPatchPair_fu_190.grp_straightLineProjectorFromLayerIJtoK_fu_1464.ap_done;
    assign module_intf_54.ap_continue = 1'b1;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_straightLineProjectorFromLayerIJtoK_fu_218.ap_start;
    assign module_intf_55.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_straightLineProjectorFromLayerIJtoK_fu_218.ap_ready;
    assign module_intf_55.ap_done = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.grp_straightLineProjectorFromLayerIJtoK_fu_218.ap_done;
    assign module_intf_55.ap_continue = 1'b1;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = 1'b0;
    assign module_intf_56.ap_ready = AESL_inst_MPSQ.grp_solveNextColumn_fu_336.tmp_getSolveNextColumnWhileConditional_fu_234.ap_ready;
    assign module_intf_56.ap_done = 1'b0;
    assign module_intf_56.ap_continue = 1'b0;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = AESL_inst_MPSQ.grp_initializeArrays_fu_354.ap_start;
    assign module_intf_57.ap_ready = AESL_inst_MPSQ.grp_initializeArrays_fu_354.ap_ready;
    assign module_intf_57.ap_done = AESL_inst_MPSQ.grp_initializeArrays_fu_354.ap_done;
    assign module_intf_57.ap_continue = 1'b1;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
